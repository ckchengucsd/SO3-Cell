.SUBCKT AOI21_X1 A1 A2 B VDD VSS ZN
MM5 ZN B VSS VSS nmos_rvt w=46.00n l=16n nfin=2
MM4 net2 A1 ZN VSS nmos_rvt w=46.00n l=16n nfin=2
MM3 net2 A2 VSS VSS nmos_rvt w=46.00n l=16n nfin=2
MM2 net6 B ZN VDD pmos_rvt w=46.00n l=16n nfin=2
MM1 net6 A1 VDD VDD pmos_rvt w=46.00n l=16n nfin=2
MM0 net6 A2 VDD VDD pmos_rvt w=46.00n l=16n nfin=2
.ENDS

.SUBCKT AOI22_X1 A1 A2 B1 B2 VDD VSS ZN
MM7 net1 B2 VSS VSS nmos_rvt w=46.00n l=16n nfin=2
MM6 ZN B1 net1 VSS nmos_rvt w=46.00n l=16n nfin=2
MM5 net0 A1 ZN VSS nmos_rvt w=46.00n l=16n nfin=2
MM4 VSS A2 net0 VSS nmos_rvt w=46.00n l=16n nfin=2
MM3 net2 B2 VDD VDD pmos_rvt w=46.00n l=16n nfin=2
MM2 VDD B1 net2 VDD pmos_rvt w=46.00n l=16n nfin=2
MM1 ZN A1 net2 VDD pmos_rvt w=46.00n l=16n nfin=2
MM0 net2 A2 ZN VDD pmos_rvt w=46.00n l=16n nfin=2
.ENDS

.SUBCKT DFFHQN_X1_SH CLK D VDD VSS QN
MM4 net10 net3 net12 VSS nmos_rvt w=46.0n l=16n nfin=2
MM5 VSS D net12 VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 VDD D net16 VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net10 net4 net16 VDD pmos_rvt w=46.0n l=16n nfin=2
MM6 VSS net10 net8 VSS nmos_rvt w=46.0n l=16n nfin=2
MM7 VDD net10 net8 VDD pmos_rvt w=46.0n l=16n nfin=2
MM10 net10 net3 net15 VDD pmos_rvt w=46.0n l=16n nfin=2
MM11 VDD net8 net15 VDD pmos_rvt w=46.0n l=16n nfin=2
MM8 VSS net8 net9 VSS nmos_rvt w=46.0n l=16n nfin=2
MM9 net10 net4 net9 VSS nmos_rvt w=46.0n l=16n nfin=2
MM13 net8 net3 net1 VDD pmos_rvt w=46.0n l=16n nfin=2
MM12 net8 net4 net1 VSS nmos_rvt w=46.0n l=16n nfin=2
MM14 net7 net1 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM15 net7 net1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM16 VSS net7 net6 VSS nmos_rvt w=46.0n l=16n nfin=2
MM17 net1 net3 net6 VSS nmos_rvt w=46.0n l=16n nfin=2
MM18 net1 net4 net14 VDD pmos_rvt w=46.0n l=16n nfin=2
MM19 VDD net7 net14 VDD pmos_rvt w=46.0n l=16n nfin=2
MM20 net3 CLK VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM23 net4 net3 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM24 QN net1 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM21 net3 CLK VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM22 net4 net3 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM25 QN net1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT FA_X1_SH A B CI CON SN VDD VSS
MM22 SN CI net081 VDD pmos_rvt w=46.0n l=16n nfin=2
MM21 net081 B net082 VDD pmos_rvt w=46.0n l=16n nfin=2
MM20 net082 A VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM15 SN CON net027 VDD pmos_rvt w=46.0n l=16n nfin=2
MM14 net027 CI VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM13 net027 B VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM12 net027 A VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM5 CON A net37 VDD pmos_rvt w=46.0n l=16n nfin=2
MM6 net37 B VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 net27 B VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 CON CI net27 VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 net27 A VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM25 SN CI net080 VSS nmos_rvt w=46.0n l=16n nfin=2
MM24 net080 B net079 VSS nmos_rvt w=46.0n l=16n nfin=2
MM23 net079 A VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM19 VSS CI net067 VSS nmos_rvt w=46.0n l=16n nfin=2
MM18 VSS B net067 VSS nmos_rvt w=46.0n l=16n nfin=2
MM17 VSS A net067 VSS nmos_rvt w=46.0n l=16n nfin=2
MM16 net067 CON SN VSS nmos_rvt w=46.0n l=16n nfin=2
MM11 VSS B net25 VSS nmos_rvt w=46.0n l=16n nfin=2
MM10 VSS B net36 VSS nmos_rvt w=46.0n l=16n nfin=2
MM9 VSS A net25 VSS nmos_rvt w=46.0n l=16n nfin=2
MM8 net36 A CON VSS nmos_rvt w=46.0n l=16n nfin=2
MM7 net25 CI CON VSS nmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT OAI21_X1 A1 A2 B VDD VSS ZN
MM5 VDD B ZN VDD pmos_rvt w=46.00n l=16n nfin=2
MM3 ZN A1 net7 VDD pmos_rvt w=46.00n l=16n nfin=2
MM4 VDD A2 net7 VDD pmos_rvt w=46.00n l=16n nfin=2
MM2 ZN B net0 VSS nmos_rvt w=46.00n l=16n nfin=2
MM0 VSS A1 net0 VSS nmos_rvt w=46.00n l=16n nfin=2
MM1 VSS A2 net0 VSS nmos_rvt w=46.00n l=16n nfin=2
.ENDS

.SUBCKT XNOR2_X1 A B VDD VSS Y
MM4 net015 A Y VSS nmos_rvt w=46.0n l=16n nfin=2
MM5 net015 B Y VSS nmos_rvt w=46.0n l=16n nfin=2
MM6 VSS net29 net015 VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 net29 A net43 VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 net43 B VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM11 net041 A VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM10 Y B net041 VDD pmos_rvt w=46.0n l=16n nfin=2
MM9 Y net29 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 net29 A VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net29 B VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT AND2_X1 A1 A2 VDD VSS Z
MM4 Z net10 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net10 A2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 net10 A1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM5 Z net10 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 net20 A2 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 net10 A1 net20 VSS nmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT AND2_X2 A1 A2 VDD VSS Z
MM4 Z net10 VDD VDD pmos_rvt w=92.0n l=16n nfin=4
MM1 net10 A2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 net10 A1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM5 Z net10 VSS VSS nmos_rvt w=92.0n l=16n nfin=4
MM3 net20 A2 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 net10 A1 net20 VSS nmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT AND3_X1 A1 A2 A3 VDD VSS Z
MM7 Z net10 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM6 net10 A3 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM5 net10 A2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM4 net10 A1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM3 Z net10 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 net30 A3 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM1 net20 A2 net30 VSS nmos_rvt w=46.0n l=16n nfin=2
MM0 net10 A1 net20 VSS nmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT AND3_X2 A1 A2 A3 VDD VSS Z
MM7 Z net10 VDD VDD pmos_rvt w=92.0n l=16n nfin=4
MM6 net10 A3 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM5 net10 A2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM4 net10 A1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM3 Z net10 VSS VSS nmos_rvt w=92.0n l=16n nfin=4
MM2 net30 A1 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM1 net20 A3 net30 VSS nmos_rvt w=46.0n l=16n nfin=2
MM0 net10 A2 net20 VSS nmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT AOI21_X2 A1 A2 B VDD VSS ZN
MM5 VSS B ZN VSS nmos_rvt w=92.00n l=16n nfin=4
MM4 ZN A1 net2 VSS nmos_rvt w=92.00n l=16n nfin=4
MM3 VSS A2 net2 VSS nmos_rvt w=92.00n l=16n nfin=4
MM2 ZN B net6 VDD pmos_rvt w=92.00n l=16n nfin=4
MM1 VDD A1 net6 VDD pmos_rvt w=92.00n l=16n nfin=4
MM0 VDD A2 net6 VDD pmos_rvt w=92.00n l=16n nfin=4
.ENDS

.SUBCKT AOI22_X2 A1 A2 B1 B2 VDD VSS ZN
MM7 net1 B2 VSS VSS nmos_rvt w=92.00n l=16n nfin=4
MM6 ZN B1 net1 VSS nmos_rvt w=92.00n l=16n nfin=4
MM5 net0 A1 ZN VSS nmos_rvt w=92.00n l=16n nfin=4
MM4 VSS A2 net0 VSS nmos_rvt w=92.00n l=16n nfin=4
MM3 net2 B2 VDD VDD pmos_rvt w=92.00n l=16n nfin=4
MM2 VDD B1 net2 VDD pmos_rvt w=92.00n l=16n nfin=4
MM1 ZN A1 net2 VDD pmos_rvt w=92.00n l=16n nfin=4
MM0 net2 A2 ZN VDD pmos_rvt w=92.00n l=16n nfin=4
.ENDS

.SUBCKT BUF_X1 I VDD VSS Z
MM3 Z in VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 in I VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM0 Z in VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 in I VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT BUF_X2 I VDD VSS Z
MM3 Z in VSS VSS nmos_rvt w=92.0n l=16n nfin=4
MM2 in I VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM0 Z in VDD VDD pmos_rvt w=92.0n l=16n nfin=4
MM1 in I VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT BUF_X4 I VDD VSS Z
MM3 Z in VSS VSS nmos_rvt w=184.0n l=16n nfin=8
MM2 in I VSS VSS nmos_rvt w=92.0n l=16n nfin=4
MM0 Z in VDD VDD pmos_rvt w=184.0n l=16n nfin=8
MM1 in I VDD VDD pmos_rvt w=92.0n l=16n nfin=4
.ENDS

.SUBCKT BUF_X8 I VDD VSS Z
MM3 Z in VSS VSS nmos_rvt w=368.0n l=16n nfin=16
MM2 in I VSS VSS nmos_rvt w=184.0n l=16n nfin=8
MM0 Z in VDD VDD pmos_rvt w=368.0n l=16n nfin=16
MM1 in I VDD VDD pmos_rvt w=184.0n l=16n nfin=8
.ENDS

.SUBCKT INV_X1 I VDD VSS ZN
MM0 ZN I VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM1 ZN I VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT INV_X2 I VDD VSS ZN
MM0 ZN I VSS VSS nmos_rvt w=92.00n l=16n nfin=4
MM1 ZN I VDD VDD pmos_rvt w=92.00n l=16n nfin=4
.ENDS

.SUBCKT INV_X4 I VDD VSS ZN
MM0 ZN I VSS VSS nmos_rvt w=184.00n l=16n nfin=8
MM1 ZN I VDD VDD pmos_rvt w=184.00n l=16n nfin=8
.ENDS

.SUBCKT INV_X8 I VDD VSS ZN
MM0 ZN I VSS VSS nmos_rvt w=368.00n l=16n nfin=16
MM1 ZN I VDD VDD pmos_rvt w=368.00n l=16n nfin=16
.ENDS

.SUBCKT MUX2_X1 I0 I1 S VDD VSS Z
MM11 Z net5 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM10 VSS I0 net6 VSS nmos_rvt w=46.0n l=16n nfin=2
MM9 net6 net2 net5 VSS nmos_rvt w=46.0n l=16n nfin=2
MM8 net5 S net4 VSS nmos_rvt w=46.0n l=16n nfin=2
MM7 VSS I1 net4 VSS nmos_rvt w=46.0n l=16n nfin=2
MM6 net2 S VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM5 Z net5 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM4 VDD I0 net11 VDD pmos_rvt w=46.0n l=16n nfin=2
MM3 net11 S net5 VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 net5 net2 net10 VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 VDD I1 net10 VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 net2 S VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NAND2_X1 A1 A2 VDD VSS ZN
MM3 net16 A2 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 ZN A1 net16 VSS nmos_rvt w=46.0n l=16n nfin=2
MM1 ZN A2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 ZN A1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NAND2_X2 A1 A2 VDD VSS ZN
MM3 net16 A2 VSS VSS nmos_rvt w=92.00n l=16n nfin=4
MM2 ZN A1 net16 VSS nmos_rvt w=92.00n l=16n nfin=4
MM1 ZN A2 VDD VDD pmos_rvt w=92.0n l=16n nfin=4
MM0 ZN A1 VDD VDD pmos_rvt w=92.0n l=16n nfin=4
.ENDS

.SUBCKT NAND3_X1 A1 A2 A3 VDD VSS ZN
MM5 net17 A3 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 net16 A2 net17 VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 ZN A1 net16 VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 ZN A3 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 ZN A2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 ZN A1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NAND3_X2 A1 A2 A3 VDD VSS ZN
MM5 net17 A3 VSS VSS nmos_rvt w=92.0n l=16n nfin=4
MM4 net16 A2 net17 VSS nmos_rvt w=92.0n l=16n nfin=4
MM3 ZN A1 net16 VSS nmos_rvt w=92.0n l=16n nfin=4
MM2 ZN A3 VDD VDD pmos_rvt w=92.0n l=16n nfin=4
MM1 ZN A2 VDD VDD pmos_rvt w=92.0n l=16n nfin=4
MM0 ZN A1 VDD VDD pmos_rvt w=92.0n l=16n nfin=4
.ENDS

.SUBCKT NAND4_X1 A1 A2 A3 A4 VDD VSS ZN
MM7 net18 A4 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM6 net17 A3 net18 VSS nmos_rvt w=46.0n l=16n nfin=2
MM5 net16 A2 net17 VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 ZN A1 net16 VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 ZN A4 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 ZN A3 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 ZN A2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 ZN A1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NAND4_X2 A1 A2 A3 A4 VDD VSS ZN
MM7 net18 A4 VSS VSS nmos_rvt w=92.0n l=16n nfin=4
MM6 net17 A3 net18 VSS nmos_rvt w=92.0n l=16n nfin=4
MM5 net16 A2 net17 VSS nmos_rvt w=92.0n l=16n nfin=4
MM4 ZN A1 net16 VSS nmos_rvt w=92.0n l=16n nfin=4
MM3 ZN A4 VDD VDD pmos_rvt w=92.0n l=16n nfin=4
MM2 ZN A3 VDD VDD pmos_rvt w=92.0n l=16n nfin=4
MM1 ZN A2 VDD VDD pmos_rvt w=92.0n l=16n nfin=4
MM0 ZN A1 VDD VDD pmos_rvt w=92.0n l=16n nfin=4
.ENDS

.SUBCKT NOR2_X1 A1 A2 VDD VSS ZN
MM3 VSS A1 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 VSS A2 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM1 net16 A1 ZN VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 VDD A2 net16 VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NOR2_X2 A1 A2 VDD VSS ZN
MM3 VSS A1 ZN VSS nmos_rvt w=92.0n l=16n nfin=4
MM2 VSS A2 ZN VSS nmos_rvt w=92.0n l=16n nfin=4
MM1 net16 A1 ZN VDD pmos_rvt w=92.0n l=16n nfin=4
MM0 VDD A2 net16 VDD pmos_rvt w=92.0n l=16n nfin=4
.ENDS

.SUBCKT NOR3_X1 A1 A2 A3 VDD VSS ZN
MM5 VSS A1 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 VSS A2 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 VSS A3 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 net20 A1 ZN VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net10 A2 net20 VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 VDD A3 net10 VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NOR3_X2 A1 A2 A3 VDD VSS ZN
MM5 VSS A1 ZN VSS nmos_rvt w=92.0n l=16n nfin=4
MM4 VSS A2 ZN VSS nmos_rvt w=92.0n l=16n nfin=4
MM3 VSS A3 ZN VSS nmos_rvt w=92.0n l=16n nfin=4
MM2 net20 A1 ZN VDD pmos_rvt w=92.0n l=16n nfin=4
MM1 net10 A2 net20 VDD pmos_rvt w=92.0n l=16n nfin=4
MM0 VDD A3 net10 VDD pmos_rvt w=92.0n l=16n nfin=4
.ENDS

.SUBCKT NOR4_X1 A1 A2 A3 A4 VDD VSS ZN
MM7 VSS A1 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM6 VSS A2 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM5 VSS A3 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 VSS A4 ZN VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 net30 A1 ZN VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 net20 A2 net30 VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net10 A3 net20 VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 VDD A4 net10 VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT NOR4_X2 A1 A2 A3 A4 VDD VSS ZN
MM7 VSS A1 ZN VSS nmos_rvt w=92.0n l=16n nfin=4
MM6 VSS A2 ZN VSS nmos_rvt w=92.0n l=16n nfin=4
MM5 VSS A3 ZN VSS nmos_rvt w=92.0n l=16n nfin=4
MM4 VSS A4 ZN VSS nmos_rvt w=92.0n l=16n nfin=4
MM3 net30 A1 ZN VDD pmos_rvt w=92.0n l=16n nfin=4
MM2 net20 A2 net30 VDD pmos_rvt w=92.0n l=16n nfin=4
MM1 net10 A3 net20 VDD pmos_rvt w=92.0n l=16n nfin=4
MM0 VDD A4 net10 VDD pmos_rvt w=92.0n l=16n nfin=4
.ENDS

.SUBCKT OAI21_X2 A1 A2 B VDD VSS ZN
MM5 VDD B ZN VDD pmos_rvt w=92.00n l=16n nfin=4
MM3 ZN A1 net7 VDD pmos_rvt w=92.00n l=16n nfin=4
MM4 VDD A2 net7 VDD pmos_rvt w=92.00n l=16n nfin=4
MM2 ZN B net0 VSS nmos_rvt w=92.00n l=16n nfin=4
MM0 VSS A1 net0 VSS nmos_rvt w=92.00n l=16n nfin=4
MM1 VSS A2 net0 VSS nmos_rvt w=92.00n l=16n nfin=4
.ENDS

.SUBCKT OAI22_X1 A1 A2 B1 B2 VDD VSS ZN
MM7 VDD B2 net8 VDD pmos_rvt w=46.00n l=16n nfin=2
MM6 ZN B1 net8 VDD pmos_rvt w=46.00n l=16n nfin=2
MM4 net9 A1 ZN VDD pmos_rvt w=46.00n l=16n nfin=2
MM5 VDD A2 net9 VDD pmos_rvt w=46.00n l=16n nfin=2
MM3 VSS B2 net2 VSS nmos_rvt w=46.00n l=16n nfin=2
MM2 VSS B1 net2 VSS nmos_rvt w=46.00n l=16n nfin=2
MM0 ZN A1 net2 VSS nmos_rvt w=46.00n l=16n nfin=2
MM1 ZN A2 net2 VSS nmos_rvt w=46.00n l=16n nfin=2
.ENDS

.SUBCKT OAI22_X2 A1 A2 B1 B2 VDD VSS ZN
MM7 VDD B2 net8 VDD pmos_rvt w=92.00n l=16n nfin=4
MM6 ZN B1 net8 VDD pmos_rvt w=92.00n l=16n nfin=4
MM4 net9 A1 ZN VDD pmos_rvt w=92.00n l=16n nfin=4
MM5 VDD A2 net9 VDD pmos_rvt w=92.00n l=16n nfin=4
MM3 VSS B2 net2 VSS nmos_rvt w=92.00n l=16n nfin=4
MM2 VSS B1 net2 VSS nmos_rvt w=92.00n l=16n nfin=4
MM0 ZN A1 net2 VSS nmos_rvt w=92.00n l=16n nfin=4
MM1 ZN A2 net2 VSS nmos_rvt w=92.00n l=16n nfin=4
.ENDS

.SUBCKT OR2_X1 A1 A2 VDD VSS Z
MM5 Z net2 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 VSS A1 net2 VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 VSS A2 net2 VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 Z net2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net2 A1 net6 VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 VDD A2 net6 VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT OR2_X2 A1 A2 VDD VSS Z
MM5 Z net2 VSS VSS nmos_rvt w=92.0n l=16n nfin=4
MM4 VSS A1 net2 VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 VSS A2 net2 VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 Z net2 VDD VDD pmos_rvt w=92.0n l=16n nfin=4
MM1 net2 A2 net6 VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 VDD A1 net6 VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT OR3_X1 A1 A2 A3 VDD VSS Z
MM7 Z net2 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM6 VSS A1 net2 VSS nmos_rvt w=46.0n l=16n nfin=2
MM5 VSS A2 net2 VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 VSS A3 net2 VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 Z net2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 net2 A1 net6 VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net7 A2 net6 VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 VDD A3 net7 VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT OR3_X2 A1 A2 A3 VDD VSS Z
MM7 Z net2 VSS VSS nmos_rvt w=92.0n l=16n nfin=4
MM6 VSS A1 net2 VSS nmos_rvt w=46.0n l=16n nfin=2
MM5 VSS A2 net2 VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 VSS A3 net2 VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 Z net2 VDD VDD pmos_rvt w=92.0n l=16n nfin=4
MM2 net2 A2 net6 VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net7 A3 net6 VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 VDD A1 net7 VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS


.SUBCKT XOR2_X1 A1 A2 VDD VSS Z
MM9 VSS A2 net5 VSS nmos_rvt w=46.0n l=16n nfin=2
MM8 net5 A1 Z VSS nmos_rvt w=46.0n l=16n nfin=2
MM7 VSS net2 Z VSS nmos_rvt w=46.0n l=16n nfin=2
MM6 VSS A1 net2 VSS nmos_rvt w=46.0n l=16n nfin=2
MM5 VSS A2 net2 VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 Z A2 net8 VDD pmos_rvt w=46.0n l=16n nfin=2
MM3 Z A1 net8 VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 VDD net2 net8 VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net2 A1 net7 VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 VDD A2 net7 VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT DFFRNQ_X1_SH D RN CK Q VDD VSS 
MM27 VSS CK ncki VSS nmos_rvt w=46.0n l=16n nfin=2
MM26 cki ncki VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM13 VDD CK ncki VDD pmos_rvt w=46.0n l=16n nfin=2
MM12 cki ncki VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM25 net10 D VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM24 net1 ncki net10 VSS nmos_rvt w=46.0n l=16n nfin=2
MM23 net15 cki net1 VSS nmos_rvt w=46.0n l=16n nfin=2
MM22 net12 net2 net15 VSS nmos_rvt w=46.0n l=16n nfin=2
MM21 VSS RN net12 VSS nmos_rvt w=46.0n l=16n nfin=2
MM20 net2 net1 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM19 net8 cki net2 VSS nmos_rvt w=46.0n l=16n nfin=2
MM18 net11 ncki net8 VSS nmos_rvt w=46.0n l=16n nfin=2
MM17 VSS net4 net11 VSS nmos_rvt w=46.0n l=16n nfin=2
MM16 net0 RN VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM15 net4 net8 net0 VSS nmos_rvt w=46.0n l=16n nfin=2
MM14 VSS net4 Q VSS nmos_rvt w=46.0n l=16n nfin=2
MM7 net9 RN VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM8 VDD net2 net9 VDD pmos_rvt w=46.0n l=16n nfin=2
MM9 net9 ncki net1 VDD pmos_rvt w=46.0n l=16n nfin=2
MM10 net1 cki net10 VDD pmos_rvt w=46.0n l=16n nfin=2
MM11 net10 D VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM6 net2 net1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM5 net8 ncki net2 VDD pmos_rvt w=46.0n l=16n nfin=2
MM4 net11 cki net8 VDD pmos_rvt w=46.0n l=16n nfin=2
MM3 VDD net4 net11 VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 net4 RN VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 VDD net8 net4 VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 VDD net4 Q VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT LHQ_X1 D E Q VDD VSS 
MM15 net4 E VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM14 net7 net4 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM13 net3 D VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM12 net5 net7 net3 VSS nmos_rvt w=46.0n l=16n nfin=2
MM11 net2 net4 net5 VSS nmos_rvt w=46.0n l=16n nfin=2
MM10 VSS net6 net2 VSS nmos_rvt w=46.0n l=16n nfin=2
MM9 net6 net5 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM8 Q net5 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM7 net4 E VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM6 net7 net4 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM5 net1 D VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM4 net5 net4 net1 VDD pmos_rvt w=46.0n l=16n nfin=2
MM3 net0 net7 net5 VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 VDD net6 net0 VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 net6 net5 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 Q net5 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT HA_X1 A B CON SN VDD VSS
MM4 net015 A SN VSS nmos_rvt w=46.0n l=16n nfin=2
MM5 net015 B SN VSS nmos_rvt w=46.0n l=16n nfin=2
MM6 VSS CON net015 VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 CON A net43 VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 net43 B VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM11 net041 A VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM10 SN B net041 VDD pmos_rvt w=46.0n l=16n nfin=2
MM9 SN CON VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 CON A VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 CON B VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT AOI222_X1_SH A1 A2 B1 B2 C1 C2 VDD VSS Y
MM6 net50 C2 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM5 Y C1 net50 VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 net51 B2 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 Y B1 net51 VSS nmos_rvt w=46.0n l=16n nfin=2
MM1 net49 A2 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM0 Y A1 net49 VSS nmos_rvt w=46.0n l=16n nfin=2
MM12 Y A2 net53 VDD pmos_rvt w=46.0n l=16n nfin=2
MM11 net53 B2 net27 VDD pmos_rvt w=46.0n l=16n nfin=2
MM10 net27 C2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM9 Y A1 net53 VDD pmos_rvt w=46.0n l=16n nfin=2
MM8 net53 B1 net27 VDD pmos_rvt w=46.0n l=16n nfin=2
MM7 net27 C1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT OAI222_X1_SH A1 A2 B1 B2 C1 C2 VDD VSS Y
MM7 net28 C2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM6 Y C1 net28 VDD pmos_rvt w=46.0n l=16n nfin=2
MM5 Y B1 net29 VDD pmos_rvt w=46.0n l=16n nfin=2
MM4 net29 B2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM3 Y A1 net30 VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 net30 A2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM13 net010 C2 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM12 net011 B2 net010 VSS nmos_rvt w=46.0n l=16n nfin=2
MM11 Y A2 net011 VSS nmos_rvt w=46.0n l=16n nfin=2
MM10 net010 C1 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM9 net011 B1 net010 VSS nmos_rvt w=46.0n l=16n nfin=2
MM8 Y A1 net011 VSS nmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT AOI211_X1 A1 A2 B C VDD VSS Y
MM20 Y C VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 Y B VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM4 Y A2 net32 VSS nmos_rvt w=46.0n l=16n nfin=2
MM5 net32 A1 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM21 net17 A2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 net17 A1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM6 net34 B net17 VDD pmos_rvt w=46.0n l=16n nfin=2
MM7 Y C net34 VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT OAI211_X1 A1 A2 B C VDD VSS Y
MM39 Y C VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM38 Y B VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM37 Y A1 net20 VDD pmos_rvt w=46.0n l=16n nfin=2
MM36 net20 A2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM41 VSS A2 net19 VSS nmos_rvt w=46.0n l=16n nfin=2
MM43 net10 C Y VSS nmos_rvt w=46.0n l=16n nfin=2
MM40 VSS A1 net19 VSS nmos_rvt w=46.0n l=16n nfin=2
MM42 net10 B net19 VSS nmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT AOI221_X1 A1 A2 B1 B2 C VDD VSS Y
MM28 Y C VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM27 net23 B2 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM26 Y B1 net23 VSS nmos_rvt w=46.0n l=16n nfin=2
MM2 Y A1 net24 VSS nmos_rvt w=46.0n l=16n nfin=2
MM0 net24 A2 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM1 s1 C s2 VDD pmos_rvt w=46.0n l=16n nfin=2
MM32 s2 B2 Y VDD pmos_rvt w=46.0n l=16n nfin=2
MM31 s1 A2 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM30 s2 B1 Y VDD pmos_rvt w=46.0n l=16n nfin=2
MM29 s1 A1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT OAI221_X1 A1 A2 B1 B2 C VDD VSS Y
MM12 VSS A2 net042 VSS nmos_rvt w=46.0n l=16n nfin=2
MM13 VSS A1 net042 VSS nmos_rvt w=46.0n l=16n nfin=2
MM11 Y B2 net044 VSS nmos_rvt w=46.0n l=16n nfin=2
MM10 Y B1 net044 VSS nmos_rvt w=46.0n l=16n nfin=2
MM14 net044 C net042 VSS nmos_rvt w=46.0n l=16n nfin=2
MM3 VDD A1 net048 VDD pmos_rvt w=46.0n l=16n nfin=2
MM2 Y B2 net047 VDD pmos_rvt w=46.0n l=16n nfin=2
MM0 net047 B1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM1 Y C VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM30 net048 A2 Y VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

.SUBCKT 2BDFFHQN_X1_SH CLK D0 D1 VDD VSS QN0 QN1
MM20 net3 CLK VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM21 net3 CLK VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM23 net4 net3 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM22 net4 net3 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM4_2 net10 net3 net12 VSS nmos_rvt w=46.0n l=16n nfin=2
MM5_2 VSS D0 net12 VSS nmos_rvt w=46.0n l=16n nfin=2
MM3_2 VDD D0 net16 VDD pmos_rvt w=46.0n l=16n nfin=2
MM1_2 net10 net4 net16 VDD pmos_rvt w=46.0n l=16n nfin=2
MM6_2 VSS net10 net8 VSS nmos_rvt w=46.0n l=16n nfin=2
MM7_2 VDD net10 net8 VDD pmos_rvt w=46.0n l=16n nfin=2
MM10_2 net10 net3 net15 VDD pmos_rvt w=46.0n l=16n nfin=2
MM11_2 VDD net8 net15 VDD pmos_rvt w=46.0n l=16n nfin=2
MM8_2 VSS net8 net9 VSS nmos_rvt w=46.0n l=16n nfin=2
MM9_2 net10 net4 net9 VSS nmos_rvt w=46.0n l=16n nfin=2
MM13_2 net8 net3 net1 VDD pmos_rvt w=46.0n l=16n nfin=2
MM12_2 net8 net4 net1 VSS nmos_rvt w=46.0n l=16n nfin=2
MM14_2 net7 net1 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM15_2 net7 net1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM16_2 VSS net7 net6 VSS nmos_rvt w=46.0n l=16n nfin=2
MM17_2 net1 net3 net6 VSS nmos_rvt w=46.0n l=16n nfin=2
MM18_2 net1 net4 net14 VDD pmos_rvt w=46.0n l=16n nfin=2
MM19_2 VDD net7 net14 VDD pmos_rvt w=46.0n l=16n nfin=2
MM24_2 QN0 net1 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM25_2 QN0 net1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM4_1 net10_1 net3 net12_1 VSS nmos_rvt w=46.0n l=16n nfin=2
MM5_1 VSS D1 net12_1 VSS nmos_rvt w=46.0n l=16n nfin=2
MM3_1 VDD D1 net16_1 VDD pmos_rvt w=46.0n l=16n nfin=2
MM1_1 net10_1 net4 net16_1 VDD pmos_rvt w=46.0n l=16n nfin=2
MM6_1 VSS net10_1 net8_1 VSS nmos_rvt w=46.0n l=16n nfin=2
MM7_1 VDD net10_1 net8_1 VDD pmos_rvt w=46.0n l=16n nfin=2
MM10_1 net10_1 net3 net15_1 VDD pmos_rvt w=46.0n l=16n nfin=2
MM11_1 VDD net8_1 net15_1 VDD pmos_rvt w=46.0n l=16n nfin=2
MM8_1 VSS net8_1 net9_1 VSS nmos_rvt w=46.0n l=16n nfin=2
MM9_1 net10_1 net4 net9_1 VSS nmos_rvt w=46.0n l=16n nfin=2
MM13_1 net8_1 net3 net1_1 VDD pmos_rvt w=46.0n l=16n nfin=2
MM12_1 net8_1 net4 net1_1 VSS nmos_rvt w=46.0n l=16n nfin=2
MM14_1 net7_1 net1_1 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM15_1 net7_1 net1_1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
MM16_1 VSS net7_1 net6_1 VSS nmos_rvt w=46.0n l=16n nfin=2
MM17_1 net1_1 net3 net6_1 VSS nmos_rvt w=46.0n l=16n nfin=2
MM18_1 net1_1 net4 net14_1 VDD pmos_rvt w=46.0n l=16n nfin=2
MM19_1 VDD net7_1 net14_1 VDD pmos_rvt w=46.0n l=16n nfin=2
MM24_1 QN1 net1_1 VSS VSS nmos_rvt w=46.0n l=16n nfin=2
MM25_1 QN1 net1_1 VDD VDD pmos_rvt w=46.0n l=16n nfin=2
.ENDS

