VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
CLEARANCEMEASURE EUCLIDEAN ;

SITE coresite_DH_P
    SIZE 0.0450 BY 0.2880 ;
    CLASS CORE ;
    SYMMETRY X Y ;
END coresite_DH_P

SITE coresite_DH_N
    SIZE 0.0450 BY 0.2880 ;
    CLASS CORE ;
    SYMMETRY X Y ;
END coresite_DH_N

SITE coresite
    SIZE 0.0450 BY 0.1440 ;
    CLASS CORE ;
    SYMMETRY X Y ;
END coresite

MACRO DFFRNQ_X1_DH
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRNQ_X1_DH 0 0 ;
  SIZE 0.4050 BY 0.2880 ;
  SYMMETRY X Y ;
  SITE coresite_DH_N ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.2590 0.1125 0.2450 ;
    END
  END D
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1150 0.0570 0.1010 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.3600 0.0910 0.3945 0.0770 ;
    END
  END Q
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2925 0.0430 0.3270 0.0290 ;
    END
  END RN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.4050 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.2700 0.4050 0.3060 ;
        RECT 0.0000 -0.0180 0.4050 0.0180 ;
    END
  END VSS
  OBS
      LAYER V0 ;
        RECT 0.2330 0.1970 0.2470 0.2110 ;
        RECT 0.2330 0.0290 0.2470 0.0430 ;
        RECT 0.1730 0.2210 0.1870 0.2350 ;
        RECT 0.1730 0.0530 0.1870 0.0670 ;
        RECT 0.1430 0.1730 0.1570 0.1870 ;
        RECT 0.1430 0.0530 0.1570 0.0670 ;
        RECT 0.1130 0.1970 0.1270 0.2110 ;
        RECT 0.1130 0.2210 0.1270 0.2350 ;
        RECT 0.1130 0.0290 0.1270 0.0430 ;
      LAYER M0 ;
        RECT 0.1455 0.2450 0.3720 0.2590 ;
        RECT 0.2355 0.2210 0.3045 0.2350 ;
        RECT 0.1680 0.2210 0.2025 0.2350 ;
        RECT 0.1080 0.2210 0.1470 0.2350 ;
        RECT 0.2130 0.1970 0.3945 0.2110 ;
        RECT 0.0330 0.1970 0.1920 0.2110 ;
        RECT 0.1905 0.1730 0.3045 0.1870 ;
        RECT 0.0105 0.1730 0.1620 0.1870 ;
        RECT 0.0780 0.1010 0.3720 0.1150 ;
        RECT 0.1455 0.0770 0.2820 0.0910 ;
        RECT 0.2355 0.0530 0.3720 0.0670 ;
        RECT 0.1350 0.0530 0.1920 0.0670 ;
        RECT 0.1905 0.0290 0.2520 0.0430 ;
        RECT 0.0105 0.0290 0.1470 0.0430 ;
      LAYER M1 ;
        RECT 0.1725 0.2400 0.1875 0.0480 ;
        RECT 0.1125 0.2400 0.1275 0.0240 ;
        RECT 0.2325 0.2160 0.2475 0.0240 ;
        RECT 0.1425 0.1920 0.1575 0.0480 ;
  END
END DFFRNQ_X1_DH

MACRO XOR2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2_X1 0 0 ;
  SIZE 0.2700 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0525 0.0960 0.0675 0.0240 ;
      LAYER M0 ;
        RECT 0.0450 0.0670 0.1245 0.0530 ;
        RECT 0.0450 0.0910 0.0795 0.0770 ;
    END
  END Z
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0180 0.0670 0.1920 0.0530 ;
      LAYER M1 ;
        RECT 0.0225 0.0960 0.0375 0.0240 ;
        RECT 0.1725 0.1200 0.1875 0.0480 ;
      LAYER M0 ;
        RECT 0.0180 0.0430 0.0570 0.0290 ;
        RECT 0.1575 0.1150 0.1920 0.1010 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.2370 0.0290 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2700 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2700 0.0180 ;
    END
  END VSS
  OBS
      LAYER V1 ;
        RECT 0.0230 0.0530 0.0370 0.0670 ;
        RECT 0.1730 0.0530 0.1870 0.0670 ;
      LAYER V0 ;
        RECT 0.0230 0.0290 0.0370 0.0430 ;
        RECT 0.1730 0.1010 0.1870 0.1150 ;
        RECT 0.2030 0.0770 0.2170 0.0910 ;
        RECT 0.2030 0.0530 0.2170 0.0670 ;
        RECT 0.0530 0.0770 0.0670 0.0910 ;
        RECT 0.0530 0.0530 0.0670 0.0670 ;
      LAYER M0 ;
        RECT 0.1905 0.0530 0.2250 0.0670 ;
        RECT 0.1230 0.0770 0.2595 0.0910 ;
        RECT 0.0105 0.1010 0.1245 0.1150 ;
      LAYER M1 ;
        RECT 0.2025 0.0960 0.2175 0.0240 ;
  END
END XOR2_X1

MACRO XNOR2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2_X1 0 0 ;
  SIZE 0.2700 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0525 0.0960 0.0675 0.0240 ;
      LAYER M0 ;
        RECT 0.0450 0.0670 0.0795 0.0530 ;
        RECT 0.0450 0.0910 0.1245 0.0770 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0180 0.1150 0.2250 0.1010 ;
      LAYER M1 ;
        RECT 0.0225 0.1200 0.0375 0.0480 ;
        RECT 0.2025 0.1200 0.2175 0.0240 ;
      LAYER M0 ;
        RECT 0.0180 0.1150 0.0570 0.1010 ;
        RECT 0.1980 0.0430 0.2370 0.0290 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1920 0.1010 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2700 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2700 0.0180 ;
    END
  END VSS
  OBS
      LAYER V1 ;
        RECT 0.0230 0.1010 0.0370 0.1150 ;
        RECT 0.2030 0.1010 0.2170 0.1150 ;
      LAYER V0 ;
        RECT 0.0530 0.0770 0.0670 0.0910 ;
        RECT 0.0530 0.0530 0.0670 0.0670 ;
        RECT 0.0230 0.1010 0.0370 0.1150 ;
        RECT 0.2030 0.0290 0.2170 0.0430 ;
        RECT 0.2330 0.0770 0.2470 0.0910 ;
        RECT 0.2330 0.0530 0.2470 0.0670 ;
      LAYER M0 ;
        RECT 0.0105 0.0290 0.1245 0.0430 ;
        RECT 0.1230 0.0530 0.2595 0.0670 ;
        RECT 0.1905 0.0770 0.2520 0.0910 ;
      LAYER M1 ;
        RECT 0.2325 0.0960 0.2475 0.0240 ;
  END
END XNOR2_X1

MACRO OR3_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3_X2 0 0 ;
  SIZE 0.2700 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0910 0.0570 0.0770 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1800 0.0910 0.2145 0.0770 ;
    END
  END Z
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.1150 0.1020 0.1010 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2700 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2700 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0530 0.2370 0.0670 ;
  END
END OR3_X2

MACRO OR3_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3_X1 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.1125 0.0290 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0910 0.1470 0.0770 ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1150 0.0570 0.1010 ;
    END
  END A1
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1800 0.1150 0.2145 0.1010 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0530 0.1920 0.0670 ;
  END
END OR3_X1

MACRO OR2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2_X2 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END A1
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0450 0.1150 0.0795 0.1010 ;
    END
  END Z
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.1150 0.2025 0.1010 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0780 0.0530 0.1695 0.0670 ;
        RECT 0.0330 0.0770 0.2145 0.0910 ;
  END
END OR2_X2

MACRO OR2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2_X1 0 0 ;
  SIZE 0.1800 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0430 0.0570 0.0290 ;
    END
  END A1
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1350 0.0430 0.1695 0.0290 ;
    END
  END Z
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.1150 0.1020 0.1010 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0555 0.0530 0.1470 0.0670 ;
        RECT 0.0105 0.0770 0.1470 0.0910 ;
  END
END OR2_X1

MACRO OAI22_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22_X2 0 0 ;
  SIZE 0.4500 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1980 0.1150 0.2520 0.1010 ;
      LAYER M1 ;
        RECT 0.2025 0.1200 0.2175 0.0480 ;
        RECT 0.2325 0.1200 0.2475 0.0480 ;
      LAYER M0 ;
        RECT 0.1455 0.0910 0.2250 0.0770 ;
        RECT 0.2250 0.0670 0.3945 0.0530 ;
    END
  END ZN
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0670 0.1020 0.0530 ;
    END
  END B2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.0670 0.1920 0.0530 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2580 0.0910 0.3270 0.0770 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.3480 0.0910 0.4170 0.0770 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.4500 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.4500 0.0180 ;
    END
  END VSS
  OBS
      LAYER V1 ;
        RECT 0.2030 0.1010 0.2170 0.1150 ;
        RECT 0.2330 0.1010 0.2470 0.1150 ;
      LAYER V0 ;
        RECT 0.2030 0.0770 0.2170 0.0910 ;
        RECT 0.2330 0.0530 0.2470 0.0670 ;
      LAYER M0 ;
        RECT 0.0555 0.0290 0.4395 0.0430 ;
        RECT 0.0105 0.1010 0.2145 0.1150 ;
        RECT 0.2355 0.1010 0.4395 0.1150 ;
  END
END OAI22_X2

MACRO OAI22_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22_X1 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0525 0.0960 0.0675 0.0240 ;
      LAYER M0 ;
        RECT 0.0450 0.0430 0.0795 0.0290 ;
        RECT 0.0450 0.0910 0.1245 0.0770 ;
    END
  END ZN
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1150 0.0570 0.1010 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1125 0.1010 ;
    END
  END A1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.1150 0.2025 0.1010 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  OBS
      LAYER V0 ;
        RECT 0.0530 0.0770 0.0670 0.0910 ;
        RECT 0.0530 0.0290 0.0670 0.0430 ;
      LAYER M0 ;
        RECT 0.0105 0.0530 0.2145 0.0670 ;
  END
END OAI22_X1

MACRO OAI222_X1_DH_P
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222_X1_DH_P 0 0 ;
  SIZE 0.1800 BY 0.2880 ;
  SYMMETRY X Y ;
  SITE coresite_DH_P ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.2640 0.1575 0.0240 ;
      LAYER M0 ;
        RECT 0.1005 0.0430 0.1620 0.0290 ;
        RECT 0.1005 0.1870 0.1620 0.1730 ;
        RECT 0.1350 0.2590 0.1695 0.2450 ;
    END
  END Y
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0430 0.0675 0.0290 ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.1150 0.1020 0.1010 ;
    END
  END C1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.1150 0.1575 0.1010 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.1870 0.0675 0.1730 ;
    END
  END B2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.2350 0.1575 0.2210 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.2590 0.1020 0.2450 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
        RECT 0.0000 0.2700 0.1800 0.3060 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VSS
  OBS
      LAYER V0 ;
        RECT 0.0230 0.0530 0.0370 0.0670 ;
        RECT 0.0230 0.2210 0.0370 0.2350 ;
        RECT 0.1430 0.0290 0.1570 0.0430 ;
        RECT 0.1430 0.2450 0.1570 0.2590 ;
        RECT 0.1430 0.1730 0.1570 0.1870 ;
      LAYER M0 ;
        RECT 0.0180 0.0530 0.1695 0.0670 ;
        RECT 0.0105 0.0770 0.1245 0.0910 ;
        RECT 0.0555 0.1970 0.1695 0.2110 ;
        RECT 0.0105 0.2210 0.0450 0.2350 ;
      LAYER M1 ;
        RECT 0.0225 0.2400 0.0375 0.0480 ;
  END
END OAI222_X1_DH_P

MACRO OAI222_X1_DH_N
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222_X1_DH_N 0 0 ;
  SIZE 0.1800 BY 0.2880 ;
  SYMMETRY X Y ;
  SITE coresite_DH_N ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0225 0.2400 0.0375 0.0720 ;
      LAYER M0 ;
        RECT 0.0180 0.0910 0.1245 0.0770 ;
        RECT 0.0105 0.2110 0.0450 0.1970 ;
        RECT 0.0180 0.2350 0.0795 0.2210 ;
    END
  END Y
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.0430 0.1020 0.0290 ;
    END
  END C1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1150 0.0570 0.1010 ;
    END
  END C2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.1150 0.1575 0.1010 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1870 0.0570 0.1730 ;
    END
  END A1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.1870 0.1575 0.1730 ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.2110 0.1125 0.1970 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
        RECT 0.0000 0.2700 0.1800 0.3060 ;
    END
  END VSS
  OBS
      LAYER V0 ;
        RECT 0.1130 0.0530 0.1270 0.0670 ;
        RECT 0.1130 0.2210 0.1270 0.2350 ;
        RECT 0.0230 0.0770 0.0370 0.0910 ;
        RECT 0.0230 0.2210 0.0370 0.2350 ;
        RECT 0.0230 0.1970 0.0370 0.2110 ;
        RECT 0.1430 0.0290 0.1570 0.0430 ;
        RECT 0.1430 0.2450 0.1570 0.2590 ;
      LAYER M0 ;
        RECT 0.1350 0.0290 0.1695 0.0430 ;
        RECT 0.0105 0.0530 0.1350 0.0670 ;
        RECT 0.1080 0.2210 0.1695 0.2350 ;
        RECT 0.0105 0.2450 0.1620 0.2590 ;
      LAYER M1 ;
        RECT 0.1125 0.2400 0.1275 0.0480 ;
        RECT 0.1425 0.2640 0.1575 0.0240 ;
  END
END OAI222_X1_DH_N

MACRO OAI221_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221_X1 0 0 ;
  SIZE 0.2700 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2025 0.0960 0.2175 0.0240 ;
      LAYER M0 ;
        RECT 0.1905 0.0430 0.2250 0.0290 ;
        RECT 0.1005 0.0910 0.2595 0.0770 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.0430 0.1575 0.0290 ;
    END
  END C
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0910 0.0675 0.0770 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1125 0.1010 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1575 0.1150 0.1920 0.1010 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.1150 0.2475 0.1010 ;
    END
  END B2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2700 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2700 0.0180 ;
    END
  END VSS
  OBS
      LAYER V0 ;
        RECT 0.2030 0.0770 0.2170 0.0910 ;
        RECT 0.2030 0.0290 0.2170 0.0430 ;
      LAYER M0 ;
        RECT 0.0105 0.0530 0.1245 0.0670 ;
        RECT 0.1455 0.0530 0.2595 0.0670 ;
  END
END OAI221_X1

MACRO OAI21_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21_X2 0 0 ;
  SIZE 0.3150 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0450 0.1150 0.1920 0.1010 ;
      LAYER M1 ;
        RECT 0.0525 0.1200 0.0675 0.0480 ;
        RECT 0.1725 0.1200 0.1875 0.0240 ;
      LAYER M0 ;
        RECT 0.0330 0.1150 0.0720 0.1010 ;
        RECT 0.1680 0.0430 0.2025 0.0290 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.1470 0.0290 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.0910 0.2820 0.0770 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1005 0.1150 0.2595 0.1010 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3150 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3150 0.0180 ;
    END
  END VSS
  OBS
      LAYER V1 ;
        RECT 0.0530 0.1010 0.0670 0.1150 ;
        RECT 0.1730 0.1010 0.1870 0.1150 ;
      LAYER V0 ;
        RECT 0.0530 0.1010 0.0670 0.1150 ;
        RECT 0.1730 0.0290 0.1870 0.0430 ;
      LAYER M0 ;
        RECT 0.0105 0.0530 0.3045 0.0670 ;
        RECT 0.0555 0.0770 0.1695 0.0910 ;
  END
END OAI21_X2

MACRO OAI21_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21_X1 0 0 ;
  SIZE 0.1800 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0430 0.0570 0.0290 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.0430 0.1575 0.0290 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0910 0.1695 0.0770 ;
    END
  END ZN
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1125 0.1010 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0530 0.1245 0.0670 ;
  END
END OAI21_X1

MACRO OAI211_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211_X1 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.0430 0.1020 0.0290 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.0430 0.1575 0.0290 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1005 0.0910 0.2145 0.0770 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1150 0.0570 0.1010 ;
    END
  END A2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.1150 0.2025 0.1010 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0530 0.1245 0.0670 ;
  END
END OAI211_X1

MACRO NOR4_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4_X2 0 0 ;
  SIZE 0.4050 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0430 0.1920 0.0290 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.0430 0.3720 0.0290 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0670 0.3945 0.0530 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1470 0.1010 ;
    END
  END A1
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2580 0.1150 0.3270 0.1010 ;
    END
  END A4
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.4050 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.4050 0.0180 ;
    END
  END VSS
  OBS
      LAYER V0 ;
        RECT 0.0230 0.1010 0.0370 0.1150 ;
        RECT 0.2030 0.1010 0.2170 0.1150 ;
        RECT 0.3530 0.1010 0.3670 0.1150 ;
      LAYER M1 ;
        RECT 0.0225 0.1200 0.0375 0.0240 ;
        RECT 0.2025 0.1200 0.2175 0.0240 ;
        RECT 0.3525 0.1200 0.3675 0.0240 ;
      LAYER M0 ;
        RECT 0.0555 0.0770 0.1695 0.0910 ;
        RECT 0.2355 0.0770 0.3495 0.0910 ;
        RECT 0.0105 0.1010 0.0450 0.1150 ;
        RECT 0.1905 0.1010 0.2250 0.1150 ;
        RECT 0.3480 0.1010 0.3945 0.1150 ;
      LAYER M2 ;
        RECT 0.0180 0.0290 0.3720 0.0430 ;
      LAYER V1 ;
        RECT 0.0230 0.0290 0.0370 0.0430 ;
        RECT 0.2030 0.0290 0.2170 0.0430 ;
        RECT 0.3530 0.0290 0.3670 0.0430 ;
  END
END NOR4_X2

MACRO NOR4_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4_X1 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0670 0.2145 0.0530 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0910 0.0570 0.0770 ;
    END
  END A1
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.0910 0.2025 0.0770 ;
    END
  END A4
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.1150 0.1020 0.1010 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
END NOR4_X1

MACRO NOR3_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3_X2 0 0 ;
  SIZE 0.3150 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0180 0.0910 0.1920 0.0770 ;
      LAYER M1 ;
        RECT 0.0225 0.0960 0.0375 0.0240 ;
        RECT 0.1725 0.0960 0.1875 0.0240 ;
      LAYER M0 ;
        RECT 0.0180 0.0430 0.0570 0.0290 ;
        RECT 0.1680 0.0430 0.2025 0.0290 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.1470 0.0290 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.0670 0.2595 0.0530 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.1150 0.2820 0.1010 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3150 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3150 0.0180 ;
    END
  END VSS
  OBS
      LAYER V1 ;
        RECT 0.0230 0.0770 0.0370 0.0910 ;
        RECT 0.1730 0.0770 0.1870 0.0910 ;
      LAYER V0 ;
        RECT 0.0230 0.0290 0.0370 0.0430 ;
        RECT 0.1730 0.0290 0.1870 0.0430 ;
      LAYER M0 ;
        RECT 0.0105 0.0770 0.3045 0.0910 ;
        RECT 0.0555 0.1010 0.1695 0.1150 ;
  END
END NOR3_X2

MACRO NOR3_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3_X1 0 0 ;
  SIZE 0.1800 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.0430 0.1020 0.0290 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0670 0.1245 0.0530 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0910 0.0570 0.0770 ;
    END
  END A1
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.1150 0.1575 0.1010 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
    END
  END VSS
END NOR3_X1

MACRO NOR2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_X2 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0430 0.1020 0.0290 ;
    END
  END A1
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.0670 0.1695 0.0530 ;
    END
  END ZN
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.1150 0.1920 0.1010 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0770 0.2145 0.0910 ;
  END
END NOR2_X2

MACRO NOR2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_X1 0 0 ;
  SIZE 0.1350 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.1125 0.0290 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0670 0.1245 0.0530 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1150 0.0570 0.1010 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1350 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1350 0.0180 ;
    END
  END VSS
END NOR2_X1

MACRO NAND4_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4_X2 0 0 ;
  SIZE 0.4050 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.1470 0.0290 ;
    END
  END A1
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2580 0.0430 0.3270 0.0290 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0910 0.3945 0.0770 ;
    END
  END ZN
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.1150 0.1920 0.1010 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.1150 0.3720 0.1010 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.4050 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.4050 0.0180 ;
    END
  END VSS
  OBS
      LAYER V0 ;
        RECT 0.0230 0.0290 0.0370 0.0430 ;
        RECT 0.2030 0.0290 0.2170 0.0430 ;
        RECT 0.3530 0.0290 0.3670 0.0430 ;
      LAYER M1 ;
        RECT 0.0225 0.1200 0.0375 0.0240 ;
        RECT 0.2025 0.1200 0.2175 0.0240 ;
        RECT 0.3525 0.1200 0.3675 0.0240 ;
      LAYER M0 ;
        RECT 0.0105 0.0290 0.0450 0.0430 ;
        RECT 0.1905 0.0290 0.2250 0.0430 ;
        RECT 0.3480 0.0290 0.3945 0.0430 ;
        RECT 0.0555 0.0530 0.1695 0.0670 ;
        RECT 0.2355 0.0530 0.3495 0.0670 ;
      LAYER M2 ;
        RECT 0.0180 0.1010 0.3720 0.1150 ;
      LAYER V1 ;
        RECT 0.0230 0.1010 0.0370 0.1150 ;
        RECT 0.2030 0.1010 0.2170 0.1150 ;
        RECT 0.3530 0.1010 0.3670 0.1150 ;
  END
END NAND4_X2

MACRO NAND4_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4_X1 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0670 0.0570 0.0530 ;
    END
  END A1
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.0670 0.2025 0.0530 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0910 0.2145 0.0770 ;
    END
  END ZN
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.1150 0.1020 0.1010 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
END NAND4_X1

MACRO NAND3_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3_X2 0 0 ;
  SIZE 0.3150 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0180 0.0670 0.1920 0.0530 ;
      LAYER M1 ;
        RECT 0.0225 0.1200 0.0375 0.0480 ;
        RECT 0.1725 0.1200 0.1875 0.0480 ;
      LAYER M0 ;
        RECT 0.0180 0.1150 0.0570 0.1010 ;
        RECT 0.1680 0.1150 0.2025 0.1010 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.0430 0.2820 0.0290 ;
    END
  END A1
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.0910 0.2595 0.0770 ;
    END
  END ZN
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1470 0.1010 ;
    END
  END A3
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3150 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3150 0.0180 ;
    END
  END VSS
  OBS
      LAYER V1 ;
        RECT 0.0230 0.0530 0.0370 0.0670 ;
        RECT 0.1730 0.0530 0.1870 0.0670 ;
      LAYER V0 ;
        RECT 0.0230 0.1010 0.0370 0.1150 ;
        RECT 0.1730 0.1010 0.1870 0.1150 ;
      LAYER M0 ;
        RECT 0.0555 0.0290 0.1695 0.0430 ;
        RECT 0.0105 0.0530 0.3045 0.0670 ;
  END
END NAND3_X2

MACRO NAND3_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3_X1 0 0 ;
  SIZE 0.1800 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.0430 0.1020 0.0290 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0670 0.0570 0.0530 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.0910 0.1695 0.0770 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.1150 0.1575 0.1010 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
    END
  END VSS
END NAND3_X1

MACRO NAND2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_X2 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0430 0.1020 0.0290 ;
    END
  END A1
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.0910 0.1695 0.0770 ;
    END
  END ZN
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.1150 0.1920 0.1010 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0530 0.2145 0.0670 ;
  END
END NAND2_X2

MACRO NAND2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_X1 0 0 ;
  SIZE 0.1350 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.1125 0.0290 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0910 0.1245 0.0770 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1150 0.0570 0.1010 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1350 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1350 0.0180 ;
    END
  END VSS
END NAND2_X1

MACRO MUX2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2_X1 0 0 ;
  SIZE 0.3150 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0430 0.1920 0.0290 ;
        RECT 0.0330 0.0910 0.1470 0.0770 ;
    END
  END S
  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.0430 0.2475 0.0290 ;
    END
  END I1
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2700 0.0910 0.3045 0.0770 ;
    END
  END Z
  PIN I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1125 0.1010 ;
    END
  END I0
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3150 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3150 0.0180 ;
    END
  END VSS
  OBS
      LAYER V0 ;
        RECT 0.1730 0.0770 0.1870 0.0910 ;
        RECT 0.1730 0.0530 0.1870 0.0670 ;
      LAYER M0 ;
        RECT 0.0105 0.0530 0.1920 0.0670 ;
        RECT 0.1680 0.0770 0.2025 0.0910 ;
        RECT 0.1455 0.1010 0.2820 0.1150 ;
      LAYER M1 ;
        RECT 0.1725 0.0960 0.1875 0.0240 ;
  END
END MUX2_X1

MACRO LHQ_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LHQ_X1 0 0 ;
  SIZE 0.4500 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.3375 0.0430 0.3720 0.0290 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0670 0.0450 0.0530 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1125 0.1010 ;
    END
  END E
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.4500 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.4500 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0330 0.0290 0.3045 0.0430 ;
        RECT 0.1005 0.0530 0.2820 0.0670 ;
        RECT 0.3030 0.0530 0.4395 0.0670 ;
        RECT 0.1005 0.0770 0.4170 0.0910 ;
        RECT 0.1455 0.1010 0.2370 0.1150 ;
        RECT 0.2580 0.1010 0.4395 0.1150 ;
  END
END LHQ_X1

MACRO INV_X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X8 0 0 ;
  SIZE 0.4050 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0430 0.3720 0.0290 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.1150 0.3495 0.1010 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.4050 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.4050 0.0180 ;
    END
  END VSS
END INV_X8

MACRO INV_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X4 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.0430 0.1695 0.0290 ;
    END
  END ZN
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.1150 0.1920 0.1010 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
END INV_X4

MACRO INV_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X2 0 0 ;
  SIZE 0.1350 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0430 0.1020 0.0290 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0450 0.1150 0.0795 0.1010 ;
    END
  END ZN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1350 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1350 0.0180 ;
    END
  END VSS
END INV_X2

MACRO INV_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X1 0 0 ;
  SIZE 0.0900 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0430 0.0795 0.0290 ;
    END
  END ZN
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1150 0.0675 0.1010 ;
    END
  END I
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.0900 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.0900 0.0180 ;
    END
  END VSS
END INV_X1

MACRO HA_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HA_X1 0 0 ;
  SIZE 0.2700 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0525 0.0960 0.0675 0.0240 ;
      LAYER M0 ;
        RECT 0.0450 0.0430 0.0795 0.0290 ;
        RECT 0.0450 0.0910 0.1245 0.0770 ;
    END
  END SN
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2325 0.0960 0.2475 0.0240 ;
      LAYER M0 ;
        RECT 0.1230 0.0430 0.2595 0.0290 ;
        RECT 0.1905 0.0910 0.2520 0.0770 ;
    END
  END CON
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0180 0.1150 0.2250 0.1010 ;
      LAYER M1 ;
        RECT 0.0225 0.1200 0.0375 0.0480 ;
        RECT 0.2025 0.1200 0.2175 0.0480 ;
      LAYER M0 ;
        RECT 0.0180 0.1150 0.0570 0.1010 ;
        RECT 0.1980 0.0670 0.2370 0.0530 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1920 0.1010 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2700 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2700 0.0180 ;
    END
  END VSS
  OBS
      LAYER V1 ;
        RECT 0.0230 0.1010 0.0370 0.1150 ;
        RECT 0.2030 0.1010 0.2170 0.1150 ;
      LAYER V0 ;
        RECT 0.0530 0.0770 0.0670 0.0910 ;
        RECT 0.0530 0.0290 0.0670 0.0430 ;
        RECT 0.2330 0.0770 0.2470 0.0910 ;
        RECT 0.2330 0.0290 0.2470 0.0430 ;
        RECT 0.0230 0.1010 0.0370 0.1150 ;
        RECT 0.2030 0.0530 0.2170 0.0670 ;
      LAYER M0 ;
        RECT 0.0105 0.0530 0.1245 0.0670 ;
  END
END HA_X1

MACRO FA_X1_DH
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FA_X1_DH 0 0 ;
  SIZE 0.3150 BY 0.2880 ;
  SYMMETRY X Y ;
  SITE coresite_DH_N ;
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2025 0.2160 0.2175 0.0240 ;
      LAYER M0 ;
        RECT 0.1680 0.0430 0.2250 0.0290 ;
        RECT 0.1455 0.2110 0.2250 0.1970 ;
    END
  END CON
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1350 0.0670 0.1695 0.0530 ;
    END
  END SN
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.0910 0.2820 0.0770 ;
    END
  END CI
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.1870 0.2820 0.1730 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.2590 0.2370 0.2450 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3150 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3150 0.0180 ;
        RECT 0.0000 0.2700 0.3150 0.3060 ;
    END
  END VSS
  OBS
      LAYER V0 ;
        RECT 0.2330 0.0530 0.2470 0.0670 ;
        RECT 0.2330 0.2210 0.2470 0.2350 ;
        RECT 0.2030 0.0290 0.2170 0.0430 ;
        RECT 0.2030 0.1970 0.2170 0.2110 ;
      LAYER M0 ;
        RECT 0.1905 0.0530 0.3045 0.0670 ;
        RECT 0.1905 0.1010 0.3045 0.1150 ;
        RECT 0.0105 0.1970 0.1245 0.2110 ;
        RECT 0.0105 0.2210 0.1245 0.2350 ;
        RECT 0.2250 0.2210 0.3045 0.2350 ;
      LAYER M1 ;
        RECT 0.2325 0.2400 0.2475 0.0480 ;
  END
END FA_X1_DH

MACRO DFFHQN_X1_DH
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQN_X1_DH 0 0 ;
  SIZE 0.3150 BY 0.2880 ;
  SYMMETRY X Y ;
  SITE coresite_DH_N ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2580 0.0430 0.2925 0.0290 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.1150 0.2475 0.1010 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.1870 0.0450 0.1730 ;
    END
  END QN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3150 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3150 0.0180 ;
        RECT 0.0000 0.2700 0.3150 0.3060 ;
    END
  END VSS
  OBS
      LAYER V0 ;
        RECT 0.1430 0.0290 0.1570 0.0430 ;
        RECT 0.1430 0.1730 0.1570 0.1870 ;
        RECT 0.2030 0.0770 0.2170 0.0910 ;
        RECT 0.2030 0.0530 0.2170 0.0670 ;
        RECT 0.2030 0.2450 0.2170 0.2590 ;
        RECT 0.0530 0.0290 0.0670 0.0430 ;
        RECT 0.0530 0.1970 0.0670 0.2110 ;
        RECT 0.1130 0.1010 0.1270 0.1150 ;
        RECT 0.1130 0.0530 0.1270 0.0670 ;
        RECT 0.1130 0.2450 0.1270 0.2590 ;
      LAYER M0 ;
        RECT 0.0450 0.0290 0.1020 0.0430 ;
        RECT 0.1350 0.0290 0.1695 0.0430 ;
        RECT 0.0105 0.0530 0.1470 0.0670 ;
        RECT 0.1680 0.0530 0.2250 0.0670 ;
        RECT 0.0330 0.0770 0.3045 0.0910 ;
        RECT 0.1080 0.1010 0.1920 0.1150 ;
        RECT 0.0780 0.1730 0.1620 0.1870 ;
        RECT 0.0450 0.1970 0.1245 0.2110 ;
        RECT 0.2130 0.1970 0.3045 0.2110 ;
        RECT 0.0330 0.2210 0.2820 0.2350 ;
        RECT 0.1080 0.2450 0.1470 0.2590 ;
        RECT 0.1680 0.2450 0.2250 0.2590 ;
      LAYER M1 ;
        RECT 0.1425 0.1920 0.1575 0.0240 ;
        RECT 0.0525 0.2160 0.0675 0.0240 ;
        RECT 0.1125 0.2640 0.1275 0.0480 ;
        RECT 0.2025 0.2640 0.2175 0.0480 ;
  END
END DFFHQN_X1_DH

MACRO BUF_X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X8 0 0 ;
  SIZE 0.5850 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0430 0.1920 0.0290 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2355 0.1150 0.5295 0.1010 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.5850 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.5850 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0555 0.0530 0.5520 0.0670 ;
  END
END BUF_X8

MACRO BUF_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X4 0 0 ;
  SIZE 0.3150 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.0430 0.2820 0.0290 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.1150 0.1695 0.1010 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3150 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3150 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0330 0.0530 0.2595 0.0670 ;
  END
END BUF_X4

MACRO BUF_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X2 0 0 ;
  SIZE 0.1800 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.0430 0.1575 0.0290 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.0910 0.0900 0.0770 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0330 0.1010 0.1695 0.1150 ;
  END
END BUF_X2

MACRO BUF_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X1 0 0 ;
  SIZE 0.1350 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0430 0.0570 0.0290 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0900 0.0910 0.1245 0.0770 ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1350 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1350 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0105 0.1010 0.1020 0.1150 ;
  END
END BUF_X1

MACRO AOI22_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22_X2 0 0 ;
  SIZE 0.4500 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1980 0.0670 0.2520 0.0530 ;
      LAYER M1 ;
        RECT 0.2025 0.0960 0.2175 0.0240 ;
        RECT 0.2325 0.1200 0.2475 0.0480 ;
      LAYER M0 ;
        RECT 0.1455 0.0430 0.2250 0.0290 ;
        RECT 0.2250 0.1150 0.3945 0.1010 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2580 0.0430 0.3270 0.0290 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.3480 0.0430 0.4170 0.0290 ;
    END
  END A2
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.1150 0.1020 0.1010 ;
    END
  END B2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.1150 0.1920 0.1010 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.4500 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.4500 0.0180 ;
    END
  END VSS
  OBS
      LAYER V1 ;
        RECT 0.2030 0.0530 0.2170 0.0670 ;
        RECT 0.2330 0.0530 0.2470 0.0670 ;
      LAYER V0 ;
        RECT 0.2030 0.0290 0.2170 0.0430 ;
        RECT 0.2330 0.1010 0.2470 0.1150 ;
      LAYER M0 ;
        RECT 0.0105 0.0530 0.2145 0.0670 ;
        RECT 0.2355 0.0530 0.4395 0.0670 ;
        RECT 0.0555 0.0770 0.4395 0.0910 ;
  END
END AOI22_X2

MACRO AOI22_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22_X1 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0525 0.1200 0.0675 0.0240 ;
      LAYER M0 ;
        RECT 0.0450 0.0430 0.1245 0.0290 ;
        RECT 0.0450 0.1150 0.0795 0.1010 ;
    END
  END ZN
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.0430 0.2025 0.0290 ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0670 0.0570 0.0530 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0670 0.1125 0.0530 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.1150 0.1470 0.1010 ;
    END
  END B1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  OBS
      LAYER V0 ;
        RECT 0.0530 0.1010 0.0670 0.1150 ;
        RECT 0.0530 0.0290 0.0670 0.0430 ;
      LAYER M0 ;
        RECT 0.0105 0.0770 0.2145 0.0910 ;
  END
END AOI22_X1

MACRO AOI222_X1_DH_P
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222_X1_DH_P 0 0 ;
  SIZE 0.1800 BY 0.2880 ;
  SYMMETRY X Y ;
  SITE coresite_DH_P ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1125 0.2160 0.1275 0.0480 ;
      LAYER M0 ;
        RECT 0.1005 0.0670 0.1350 0.0530 ;
        RECT 0.1080 0.1150 0.1695 0.1010 ;
        RECT 0.0555 0.2110 0.1350 0.1970 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.0910 0.1020 0.0770 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.0910 0.1575 0.0770 ;
    END
  END A1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1150 0.0570 0.1010 ;
    END
  END B2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1870 0.0570 0.1730 ;
    END
  END B1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.1870 0.1575 0.1730 ;
    END
  END C2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.2590 0.1125 0.2450 ;
    END
  END C1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
        RECT 0.0000 0.2700 0.1800 0.3060 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VSS
  OBS
      LAYER V0 ;
        RECT 0.1130 0.1010 0.1270 0.1150 ;
        RECT 0.1130 0.0530 0.1270 0.0670 ;
        RECT 0.1130 0.1970 0.1270 0.2110 ;
        RECT 0.0530 0.0530 0.0670 0.0670 ;
        RECT 0.0530 0.2210 0.0670 0.2350 ;
        RECT 0.0230 0.0290 0.0370 0.0430 ;
        RECT 0.0230 0.2450 0.0370 0.2590 ;
      LAYER M0 ;
        RECT 0.0180 0.0290 0.1695 0.0430 ;
        RECT 0.0105 0.0530 0.0720 0.0670 ;
        RECT 0.0450 0.2210 0.1695 0.2350 ;
        RECT 0.0105 0.2450 0.0450 0.2590 ;
      LAYER M1 ;
        RECT 0.0525 0.2400 0.0675 0.0480 ;
        RECT 0.0225 0.2640 0.0375 0.0240 ;
  END
END AOI222_X1_DH_P

MACRO AOI222_X1_DH_N
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222_X1_DH_N 0 0 ;
  SIZE 0.1800 BY 0.2880 ;
  SYMMETRY X Y ;
  SITE coresite_DH_N ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.1425 0.2640 0.1575 0.0240 ;
      LAYER M0 ;
        RECT 0.1350 0.0430 0.1695 0.0290 ;
        RECT 0.1005 0.1150 0.1620 0.1010 ;
        RECT 0.1005 0.2590 0.1620 0.2450 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.0430 0.1020 0.0290 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.0670 0.1575 0.0530 ;
    END
  END A1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1150 0.0570 0.1010 ;
    END
  END B2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.1870 0.1020 0.1730 ;
    END
  END C1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.1870 0.1575 0.1730 ;
    END
  END B1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.2590 0.0570 0.2450 ;
    END
  END C2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
        RECT 0.0000 0.2700 0.1800 0.3060 ;
    END
  END VSS
  OBS
      LAYER V0 ;
        RECT 0.1430 0.1010 0.1570 0.1150 ;
        RECT 0.1430 0.0290 0.1570 0.0430 ;
        RECT 0.1430 0.2450 0.1570 0.2590 ;
        RECT 0.0230 0.0530 0.0370 0.0670 ;
        RECT 0.0230 0.2210 0.0370 0.2350 ;
      LAYER M0 ;
        RECT 0.0105 0.0530 0.0450 0.0670 ;
        RECT 0.0555 0.0770 0.1695 0.0910 ;
        RECT 0.0105 0.1970 0.1245 0.2110 ;
        RECT 0.0180 0.2210 0.1695 0.2350 ;
      LAYER M1 ;
        RECT 0.0225 0.2400 0.0375 0.0480 ;
  END
END AOI222_X1_DH_N

MACRO AOI221_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221_X1 0 0 ;
  SIZE 0.2700 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0525 0.1200 0.0675 0.0480 ;
      LAYER M0 ;
        RECT 0.0105 0.0670 0.1695 0.0530 ;
        RECT 0.0450 0.1150 0.0795 0.1010 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0430 0.0570 0.0290 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.1125 0.0290 ;
    END
  END B2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1575 0.0430 0.1920 0.0290 ;
    END
  END A1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.1150 0.1470 0.1010 ;
    END
  END C
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.1150 0.2475 0.1010 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2700 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2700 0.0180 ;
    END
  END VSS
  OBS
      LAYER V0 ;
        RECT 0.0530 0.1010 0.0670 0.1150 ;
        RECT 0.0530 0.0530 0.0670 0.0670 ;
      LAYER M0 ;
        RECT 0.0105 0.0770 0.1245 0.0910 ;
        RECT 0.1455 0.0770 0.2595 0.0910 ;
  END
END AOI221_X1

MACRO AOI21_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21_X2 0 0 ;
  SIZE 0.3150 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0450 0.0670 0.1920 0.0530 ;
      LAYER M1 ;
        RECT 0.0525 0.0960 0.0675 0.0240 ;
        RECT 0.1725 0.1200 0.1875 0.0480 ;
      LAYER M0 ;
        RECT 0.0330 0.0430 0.0720 0.0290 ;
        RECT 0.1680 0.1150 0.2025 0.1010 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1005 0.0430 0.2595 0.0290 ;
    END
  END ZN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.0670 0.2820 0.0530 ;
    END
  END B
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1470 0.1010 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3150 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3150 0.0180 ;
    END
  END VSS
  OBS
      LAYER V1 ;
        RECT 0.0530 0.0530 0.0670 0.0670 ;
        RECT 0.1730 0.0530 0.1870 0.0670 ;
      LAYER V0 ;
        RECT 0.0530 0.0290 0.0670 0.0430 ;
        RECT 0.1730 0.1010 0.1870 0.1150 ;
      LAYER M0 ;
        RECT 0.0555 0.0530 0.1695 0.0670 ;
        RECT 0.0105 0.0770 0.3045 0.0910 ;
  END
END AOI21_X2

MACRO AOI21_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21_X1 0 0 ;
  SIZE 0.1800 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0430 0.0570 0.0290 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.0430 0.1575 0.0290 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0670 0.1695 0.0530 ;
    END
  END ZN
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.1150 0.1020 0.1010 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0770 0.1245 0.0910 ;
  END
END AOI21_X1

MACRO AOI211_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211_X1 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0430 0.0570 0.0290 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1005 0.0670 0.2145 0.0530 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1125 0.1010 ;
    END
  END A2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.1150 0.2025 0.1010 ;
    END
  END C
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0770 0.1245 0.0910 ;
  END
END AOI211_X1

MACRO AND3_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3_X2 0 0 ;
  SIZE 0.2700 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.0430 0.2025 0.0290 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.0670 0.0900 0.0530 ;
    END
  END Z
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.0670 0.2475 0.0530 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.1150 0.1470 0.1010 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2700 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2700 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0330 0.0770 0.2595 0.0910 ;
  END
END AND3_X2

MACRO AND3_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3_X1 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0670 0.0570 0.0530 ;
    END
  END A1
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1800 0.0670 0.2145 0.0530 ;
    END
  END Z
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1125 0.1010 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0770 0.1920 0.0910 ;
  END
END AND3_X1

MACRO AND2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_X2 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0450 0.1150 0.0795 0.1010 ;
    END
  END Z
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.1150 0.2025 0.1010 ;
    END
  END A1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0330 0.0530 0.2145 0.0670 ;
        RECT 0.0780 0.0770 0.1695 0.0910 ;
  END
END AND2_X2

MACRO AND2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_X1 0 0 ;
  SIZE 0.1800 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0430 0.0570 0.0290 ;
    END
  END A1
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1350 0.0430 0.1695 0.0290 ;
    END
  END Z
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.1150 0.1020 0.1010 ;
    END
  END A2
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
    END
  END VSS
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0530 0.1470 0.0670 ;
        RECT 0.0555 0.0770 0.1470 0.0910 ;
  END
END AND2_X1

MACRO 2BDFFHQN_X1_DH
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN 2BDFFHQN_X1_DH 0 0 ;
  SIZE 0.5850 BY 0.2880 ;
  SYMMETRY X Y ;
  SITE coresite_DH_N ;
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.4725 0.2590 0.5070 0.2450 ;
    END
  END D0
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.2350 0.0450 0.2210 ;
    END
  END QN0
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.5280 0.0670 0.5625 0.0530 ;
    END
  END CLK
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.4725 0.0910 0.5070 0.0770 ;
    END
  END D1
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0430 0.0450 0.0290 ;
    END
  END QN1
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.5850 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.2700 0.5850 0.3060 ;
        RECT 0.0000 -0.0180 0.5850 0.0180 ;
    END
  END VSS
  OBS
      LAYER V0 ;
        RECT 0.3830 0.1730 0.3970 0.1870 ;
        RECT 0.3830 0.2210 0.3970 0.2350 ;
        RECT 0.3830 0.0290 0.3970 0.0430 ;
        RECT 0.2330 0.2450 0.2470 0.2590 ;
        RECT 0.2330 0.0530 0.2470 0.0670 ;
        RECT 0.2330 0.1010 0.2470 0.1150 ;
      LAYER M0 ;
        RECT 0.3030 0.2450 0.4395 0.2590 ;
        RECT 0.2130 0.2450 0.2520 0.2590 ;
        RECT 0.1005 0.2450 0.1920 0.2590 ;
        RECT 0.4380 0.2210 0.5520 0.2350 ;
        RECT 0.2580 0.2210 0.4170 0.2350 ;
        RECT 0.3930 0.1970 0.5520 0.2110 ;
        RECT 0.2805 0.1970 0.3720 0.2110 ;
        RECT 0.0330 0.1970 0.2595 0.2110 ;
        RECT 0.2130 0.1730 0.5745 0.1870 ;
        RECT 0.2280 0.1010 0.5745 0.1150 ;
        RECT 0.2805 0.0770 0.3720 0.0910 ;
        RECT 0.0330 0.0770 0.2595 0.0910 ;
        RECT 0.3030 0.0530 0.4395 0.0670 ;
        RECT 0.2130 0.0530 0.2520 0.0670 ;
        RECT 0.1005 0.0530 0.1920 0.0670 ;
        RECT 0.4380 0.0290 0.5745 0.0430 ;
        RECT 0.2580 0.0290 0.4170 0.0430 ;
      LAYER M1 ;
        RECT 0.2325 0.2640 0.2475 0.0480 ;
        RECT 0.3825 0.2400 0.3975 0.0240 ;
  END
END 2BDFFHQN_X1_DH

MACRO AOI222_X1_SH
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222_X1_SH 0 0 ;
  SIZE 0.3600 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.0430 0.2025 0.0290 ;
    END
  END B2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2475 0.0430 0.2820 0.0290 ;
    END
  END A1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0670 0.0570 0.0530 ;
    END
  END C2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1005 0.0670 0.2595 0.0530 ;
        RECT 0.2355 0.0910 0.3495 0.0770 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.3030 0.0670 0.3375 0.0530 ;
    END
  END A2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1125 0.1010 ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3600 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3600 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0770 0.2145 0.0910 ;
        RECT 0.1455 0.1010 0.3045 0.1150 ;
  END
END AOI222_X1_SH

MACRO OAI222_X1_SH
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222_X1_SH 0 0 ;
  SIZE 0.3600 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.1125 0.0290 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2355 0.0670 0.3495 0.0530 ;
        RECT 0.1005 0.0910 0.2595 0.0770 ;
    END
  END Y
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0910 0.0570 0.0770 ;
    END
  END C2
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.3030 0.0910 0.3375 0.0770 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.1150 0.1470 0.1010 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.1150 0.2025 0.1010 ;
    END
  END B2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2475 0.1150 0.2820 0.1010 ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3600 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3600 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.1455 0.0290 0.3045 0.0430 ;
        RECT 0.0105 0.0530 0.2145 0.0670 ;
  END
END OAI222_X1_SH
