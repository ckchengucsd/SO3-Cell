VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
CLEARANCEMEASURE EUCLIDEAN ;

SITE coresite
    SIZE 0.0450 BY 0.1440 ;
    CLASS CORE ;
    SYMMETRY Y ;
END coresite

MACRO XNOR2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2_X1 0 0 ;
  SIZE 0.2700 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0525 0.0960 0.0675 0.0240 ;
      LAYER M0 ;
        RECT 0.0450 0.0670 0.0795 0.0530 ;
        RECT 0.0450 0.0910 0.1245 0.0770 ;
    END
  END Y
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0180 0.1150 0.2250 0.1010 ;
      LAYER M1 ;
        RECT 0.0225 0.1200 0.0375 0.0480 ;
        RECT 0.2025 0.1200 0.2175 0.0240 ;
      LAYER M0 ;
        RECT 0.0180 0.1150 0.0570 0.1010 ;
        RECT 0.1980 0.0430 0.2370 0.0290 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1920 0.1010 ;
    END
  END B
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2700 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2700 0.1620 ;
    END
  END VDD
  OBS
      LAYER V1 ;
        RECT 0.0230 0.1010 0.0370 0.1150 ;
        RECT 0.2030 0.1010 0.2170 0.1150 ;
      LAYER M0 ;
        RECT 0.0105 0.0290 0.1245 0.0430 ;
        RECT 0.1230 0.0530 0.2595 0.0670 ;
        RECT 0.1905 0.0770 0.2520 0.0910 ;
      LAYER V0 ;
        RECT 0.0530 0.0770 0.0670 0.0910 ;
        RECT 0.0530 0.0530 0.0670 0.0670 ;
        RECT 0.0230 0.1010 0.0370 0.1150 ;
        RECT 0.2030 0.0290 0.2170 0.0430 ;
        RECT 0.2330 0.0770 0.2470 0.0910 ;
        RECT 0.2330 0.0530 0.2470 0.0670 ;
      LAYER M1 ;
        RECT 0.2325 0.0960 0.2475 0.0240 ;
  END
END XNOR2_X1

MACRO OAI222_X1_SH
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI222_X1_SH 0 0 ;
  SIZE 0.3600 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.1125 0.0290 ;
    END
  END C1
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2355 0.0670 0.3495 0.0530 ;
        RECT 0.1005 0.0910 0.2595 0.0770 ;
    END
  END Y
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0910 0.0570 0.0770 ;
    END
  END C2
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.3030 0.0910 0.3375 0.0770 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.1150 0.1470 0.1010 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.1150 0.2025 0.1010 ;
    END
  END B2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2475 0.1150 0.2820 0.1010 ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3600 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3600 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.1455 0.0290 0.3045 0.0430 ;
        RECT 0.0105 0.0530 0.2145 0.0670 ;
  END
END OAI222_X1_SH

MACRO OAI221_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI221_X1 0 0 ;
  SIZE 0.2700 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2025 0.0960 0.2175 0.0240 ;
      LAYER M0 ;
        RECT 0.1905 0.0430 0.2250 0.0290 ;
        RECT 0.1005 0.0910 0.2595 0.0770 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.0430 0.1575 0.0290 ;
    END
  END C
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0910 0.0675 0.0770 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1125 0.1010 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1575 0.1150 0.1920 0.1010 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.1150 0.2475 0.1010 ;
    END
  END B2
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2700 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2700 0.1620 ;
    END
  END VDD
  OBS
      LAYER V0 ;
        RECT 0.2030 0.0770 0.2170 0.0910 ;
        RECT 0.2030 0.0290 0.2170 0.0430 ;
      LAYER M0 ;
        RECT 0.0105 0.0530 0.1245 0.0670 ;
        RECT 0.1455 0.0530 0.2595 0.0670 ;
  END
END OAI221_X1

MACRO OAI211_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI211_X1 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.0430 0.1020 0.0290 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.0430 0.1575 0.0290 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1005 0.0910 0.2145 0.0770 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1150 0.0570 0.1010 ;
    END
  END A2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.1150 0.2025 0.1010 ;
    END
  END C
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0530 0.1245 0.0670 ;
  END
END OAI211_X1

MACRO HA_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN HA_X1 0 0 ;
  SIZE 0.2700 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0525 0.0960 0.0675 0.0240 ;
      LAYER M0 ;
        RECT 0.0450 0.0430 0.0795 0.0290 ;
        RECT 0.0450 0.0910 0.1245 0.0770 ;
    END
  END SN
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.2325 0.0960 0.2475 0.0240 ;
      LAYER M0 ;
        RECT 0.1230 0.0430 0.2595 0.0290 ;
        RECT 0.1905 0.0910 0.2520 0.0770 ;
    END
  END CON
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0180 0.1150 0.2250 0.1010 ;
      LAYER M1 ;
        RECT 0.0225 0.1200 0.0375 0.0480 ;
        RECT 0.2025 0.1200 0.2175 0.0480 ;
      LAYER M0 ;
        RECT 0.0180 0.1150 0.0570 0.1010 ;
        RECT 0.1980 0.0670 0.2370 0.0530 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1920 0.1010 ;
    END
  END B
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2700 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2700 0.1620 ;
    END
  END VDD
  OBS
      LAYER V1 ;
        RECT 0.0230 0.1010 0.0370 0.1150 ;
        RECT 0.2030 0.1010 0.2170 0.1150 ;
      LAYER V0 ;
        RECT 0.0530 0.0770 0.0670 0.0910 ;
        RECT 0.0530 0.0290 0.0670 0.0430 ;
        RECT 0.2330 0.0770 0.2470 0.0910 ;
        RECT 0.2330 0.0290 0.2470 0.0430 ;
        RECT 0.0230 0.1010 0.0370 0.1150 ;
        RECT 0.2030 0.0530 0.2170 0.0670 ;
      LAYER M0 ;
        RECT 0.0105 0.0530 0.1245 0.0670 ;
  END
END HA_X1

MACRO FA_X1_SH
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FA_X1_SH 0 0 ;
  SIZE 0.5850 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0450 0.0910 0.4950 0.0770 ;
      LAYER M1 ;
        RECT 0.2025 0.0960 0.2175 0.0240 ;
        RECT 0.4725 0.0960 0.4875 0.0240 ;
        RECT 0.0525 0.1200 0.0675 0.0480 ;
      LAYER M0 ;
        RECT 0.1680 0.0910 0.2820 0.0770 ;
        RECT 0.4680 0.0430 0.5070 0.0290 ;
        RECT 0.0330 0.1150 0.0720 0.1010 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3150 0.1150 0.5220 0.1010 ;
      LAYER M1 ;
        RECT 0.3225 0.1200 0.3375 0.0480 ;
        RECT 0.5025 0.1200 0.5175 0.0480 ;
      LAYER M0 ;
        RECT 0.0780 0.0670 0.3420 0.0530 ;
        RECT 0.4950 0.1150 0.5520 0.1010 ;
    END
  END B
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1455 0.0430 0.4170 0.0290 ;
    END
  END CON
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.3600 0.0910 0.3945 0.0770 ;
    END
  END SN
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.1150 0.4620 0.1010 ;
    END
  END CI
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.5850 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.5850 0.1620 ;
    END
  END VDD
  OBS
      LAYER V1 ;
        RECT 0.0530 0.0770 0.0670 0.0910 ;
        RECT 0.2030 0.0770 0.2170 0.0910 ;
        RECT 0.4730 0.0770 0.4870 0.0910 ;
        RECT 0.3230 0.1010 0.3370 0.1150 ;
        RECT 0.5030 0.1010 0.5170 0.1150 ;
      LAYER V0 ;
        RECT 0.0530 0.1010 0.0670 0.1150 ;
        RECT 0.2030 0.0770 0.2170 0.0910 ;
        RECT 0.4730 0.0290 0.4870 0.0430 ;
        RECT 0.3230 0.0530 0.3370 0.0670 ;
        RECT 0.5030 0.1010 0.5170 0.1150 ;
      LAYER M0 ;
        RECT 0.0105 0.0290 0.1245 0.0430 ;
        RECT 0.4155 0.0530 0.5295 0.0670 ;
        RECT 0.0105 0.0770 0.1245 0.0910 ;
        RECT 0.4155 0.0770 0.5295 0.0910 ;
  END
END FA_X1_SH

MACRO AOI222_X1_SH
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI222_X1_SH 0 0 ;
  SIZE 0.3600 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.0430 0.2025 0.0290 ;
    END
  END B2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2475 0.0430 0.2820 0.0290 ;
    END
  END A1
  PIN C2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0670 0.0570 0.0530 ;
    END
  END C2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1005 0.0670 0.2595 0.0530 ;
        RECT 0.2355 0.0910 0.3495 0.0770 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.3030 0.0670 0.3375 0.0530 ;
    END
  END A2
  PIN C1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1125 0.1010 ;
    END
  END C1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3600 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3600 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0770 0.2145 0.0910 ;
        RECT 0.1455 0.1010 0.3045 0.1150 ;
  END
END AOI222_X1_SH

MACRO AOI221_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI221_X1 0 0 ;
  SIZE 0.2700 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0525 0.1200 0.0675 0.0480 ;
      LAYER M0 ;
        RECT 0.0105 0.0670 0.1695 0.0530 ;
        RECT 0.0450 0.1150 0.0795 0.1010 ;
    END
  END Y
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0430 0.0570 0.0290 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.1125 0.0290 ;
    END
  END B2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1575 0.0430 0.1920 0.0290 ;
    END
  END A1
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.1150 0.1470 0.1010 ;
    END
  END C
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.1150 0.2475 0.1010 ;
    END
  END A2
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2700 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2700 0.1620 ;
    END
  END VDD
  OBS
      LAYER V0 ;
        RECT 0.0530 0.1010 0.0670 0.1150 ;
        RECT 0.0530 0.0530 0.0670 0.0670 ;
      LAYER M0 ;
        RECT 0.0105 0.0770 0.1245 0.0910 ;
        RECT 0.1455 0.0770 0.2595 0.0910 ;
  END
END AOI221_X1

MACRO AOI211_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI211_X1 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0430 0.0570 0.0290 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1005 0.0670 0.2145 0.0530 ;
    END
  END Y
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1125 0.1010 ;
    END
  END A2
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.1150 0.2025 0.1010 ;
    END
  END C
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0770 0.1245 0.0910 ;
  END
END AOI211_X1

MACRO 2BDFFHQN_X1_SH
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN 2BDFFHQN_X1_SH 0 0 ;
  SIZE 1.1250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN QN0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 1.0005 0.0910 1.0350 0.0770 ;
    END
  END QN0
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.5730 0.0910 0.6075 0.0770 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.5175 0.0910 0.5520 0.0770 ;
    END
  END D1
  PIN QN1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0910 0.0450 0.0770 ;
    END
  END QN1
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 1.0680 0.0670 1.1025 0.0530 ;
    END
  END CLK
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 1.1250 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 1.1250 0.0180 ;
    END
  END VSS
  OBS
      LAYER M2 ;
        RECT 0.6480 0.0770 0.7020 0.0910 ;
        RECT 0.2880 0.0770 0.3420 0.0910 ;
      LAYER V0 ;
        RECT 0.6830 0.1010 0.6970 0.1150 ;
        RECT 0.6530 0.0530 0.6670 0.0670 ;
        RECT 0.4430 0.0530 0.4570 0.0670 ;
        RECT 0.4430 0.1010 0.4570 0.1150 ;
        RECT 0.2630 0.0290 0.2770 0.0430 ;
        RECT 0.2630 0.1010 0.2770 0.1150 ;
        RECT 0.8030 0.0290 0.8170 0.0430 ;
        RECT 0.8030 0.0770 0.8170 0.0910 ;
        RECT 0.5630 0.0290 0.5770 0.0430 ;
        RECT 0.5630 0.1010 0.5770 0.1150 ;
        RECT 0.3230 0.0290 0.3370 0.0430 ;
        RECT 0.2930 0.0770 0.3070 0.0910 ;
      LAYER M1 ;
        RECT 0.6825 0.1200 0.6975 0.0480 ;
        RECT 0.5625 0.1200 0.5775 0.0240 ;
        RECT 0.4425 0.1200 0.4575 0.0480 ;
        RECT 0.2625 0.1200 0.2775 0.0240 ;
        RECT 0.8025 0.0960 0.8175 0.0240 ;
        RECT 0.6525 0.0960 0.6675 0.0240 ;
        RECT 0.3225 0.0960 0.3375 0.0240 ;
        RECT 0.2925 0.0960 0.3075 0.0240 ;
      LAYER V1 ;
        RECT 0.6830 0.0770 0.6970 0.0910 ;
        RECT 0.6530 0.0770 0.6670 0.0910 ;
        RECT 0.3230 0.0770 0.3370 0.0910 ;
        RECT 0.2930 0.0770 0.3070 0.0910 ;
      LAYER M0 ;
        RECT 0.6630 0.1010 1.1145 0.1150 ;
        RECT 0.4830 0.1010 0.6420 0.1150 ;
        RECT 0.2580 0.1010 0.4620 0.1150 ;
        RECT 0.1005 0.1010 0.2370 0.1150 ;
        RECT 0.8880 0.0770 0.9795 0.0910 ;
        RECT 0.7980 0.0770 0.8670 0.0910 ;
        RECT 0.6405 0.0770 0.7770 0.0910 ;
        RECT 0.3480 0.0770 0.4845 0.0910 ;
        RECT 0.1455 0.0770 0.3150 0.0910 ;
        RECT 0.8205 0.0530 1.0470 0.0670 ;
        RECT 0.7080 0.0530 0.7995 0.0670 ;
        RECT 0.4380 0.0530 0.6750 0.0670 ;
        RECT 0.3255 0.0530 0.4170 0.0670 ;
        RECT 0.0330 0.0530 0.3045 0.0670 ;
        RECT 0.8430 0.0290 1.1145 0.0430 ;
        RECT 0.3030 0.0290 0.8220 0.0430 ;
        RECT 0.1680 0.0290 0.2820 0.0430 ;
  END
END 2BDFFHQN_X1_SH

MACRO XOR2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2_X1 0 0 ;
  SIZE 0.2700 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0525 0.0960 0.0675 0.0240 ;
      LAYER M0 ;
        RECT 0.0450 0.0670 0.1245 0.0530 ;
        RECT 0.0450 0.0910 0.0795 0.0770 ;
    END
  END Z
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0180 0.0670 0.1920 0.0530 ;
      LAYER M1 ;
        RECT 0.0225 0.0960 0.0375 0.0240 ;
        RECT 0.1725 0.1200 0.1875 0.0480 ;
      LAYER M0 ;
        RECT 0.0180 0.0430 0.0570 0.0290 ;
        RECT 0.1575 0.1150 0.1920 0.1010 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.2370 0.0290 ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2700 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2700 0.1620 ;
    END
  END VDD
  OBS
      LAYER V1 ;
        RECT 0.0230 0.0530 0.0370 0.0670 ;
        RECT 0.1730 0.0530 0.1870 0.0670 ;
      LAYER M0 ;
        RECT 0.1905 0.0530 0.2250 0.0670 ;
        RECT 0.1230 0.0770 0.2595 0.0910 ;
        RECT 0.0105 0.1010 0.1245 0.1150 ;
      LAYER V0 ;
        RECT 0.0230 0.0290 0.0370 0.0430 ;
        RECT 0.1730 0.1010 0.1870 0.1150 ;
        RECT 0.2030 0.0770 0.2170 0.0910 ;
        RECT 0.2030 0.0530 0.2170 0.0670 ;
        RECT 0.0530 0.0770 0.0670 0.0910 ;
        RECT 0.0530 0.0530 0.0670 0.0670 ;
      LAYER M1 ;
        RECT 0.2025 0.0960 0.2175 0.0240 ;
  END
END XOR2_X1

MACRO OR3_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3_X2 0 0 ;
  SIZE 0.2700 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0910 0.0570 0.0770 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1800 0.0910 0.2145 0.0770 ;
    END
  END Z
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.1150 0.1020 0.1010 ;
    END
  END A3
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2700 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2700 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0530 0.2370 0.0670 ;
  END
END OR3_X2

MACRO OR3_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3_X1 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.1125 0.0290 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0910 0.1470 0.0770 ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1150 0.0570 0.1010 ;
    END
  END A1
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1800 0.1150 0.2145 0.1010 ;
    END
  END Z
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0530 0.1920 0.0670 ;
  END
END OR3_X1

MACRO OR2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2_X2 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END A1
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0450 0.1150 0.0795 0.1010 ;
    END
  END Z
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.1150 0.2025 0.1010 ;
    END
  END A2
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0780 0.0530 0.1695 0.0670 ;
        RECT 0.0330 0.0770 0.2145 0.0910 ;
  END
END OR2_X2

MACRO OR2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2_X1 0 0 ;
  SIZE 0.1800 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0430 0.0570 0.0290 ;
    END
  END A1
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1350 0.0430 0.1695 0.0290 ;
    END
  END Z
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.1150 0.1020 0.1010 ;
    END
  END A2
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0555 0.0530 0.1470 0.0670 ;
        RECT 0.0105 0.0770 0.1470 0.0910 ;
  END
END OR2_X1

MACRO OAI22_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22_X2 0 0 ;
  SIZE 0.4500 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1980 0.1150 0.2520 0.1010 ;
      LAYER M1 ;
        RECT 0.2025 0.1200 0.2175 0.0480 ;
        RECT 0.2325 0.1200 0.2475 0.0480 ;
      LAYER M0 ;
        RECT 0.1455 0.0910 0.2250 0.0770 ;
        RECT 0.2250 0.0670 0.3945 0.0530 ;
    END
  END ZN
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0670 0.1020 0.0530 ;
    END
  END B2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.0670 0.1920 0.0530 ;
    END
  END B1
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2580 0.0910 0.3270 0.0770 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.3480 0.0910 0.4170 0.0770 ;
    END
  END A2
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.4500 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.4500 0.1620 ;
    END
  END VDD
  OBS
      LAYER V1 ;
        RECT 0.2030 0.1010 0.2170 0.1150 ;
        RECT 0.2330 0.1010 0.2470 0.1150 ;
      LAYER V0 ;
        RECT 0.2030 0.0770 0.2170 0.0910 ;
        RECT 0.2330 0.0530 0.2470 0.0670 ;
      LAYER M0 ;
        RECT 0.0555 0.0290 0.4395 0.0430 ;
        RECT 0.0105 0.1010 0.2145 0.1150 ;
        RECT 0.2355 0.1010 0.4395 0.1150 ;
  END
END OAI22_X2

MACRO OAI22_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22_X1 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0525 0.0960 0.0675 0.0240 ;
      LAYER M0 ;
        RECT 0.0450 0.0430 0.0795 0.0290 ;
        RECT 0.0450 0.0910 0.1245 0.0770 ;
    END
  END ZN
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END B1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1150 0.0570 0.1010 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1125 0.1010 ;
    END
  END A1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.1150 0.2025 0.1010 ;
    END
  END B2
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  OBS
      LAYER V0 ;
        RECT 0.0530 0.0770 0.0670 0.0910 ;
        RECT 0.0530 0.0290 0.0670 0.0430 ;
      LAYER M0 ;
        RECT 0.0105 0.0530 0.2145 0.0670 ;
  END
END OAI22_X1

MACRO OAI21_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21_X2 0 0 ;
  SIZE 0.3150 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0450 0.1150 0.1920 0.1010 ;
      LAYER M1 ;
        RECT 0.0525 0.1200 0.0675 0.0480 ;
        RECT 0.1725 0.1200 0.1875 0.0240 ;
      LAYER M0 ;
        RECT 0.0330 0.1150 0.0720 0.1010 ;
        RECT 0.1680 0.0430 0.2025 0.0290 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.1470 0.0290 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.0910 0.2820 0.0770 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1005 0.1150 0.2595 0.1010 ;
    END
  END ZN
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3150 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3150 0.1620 ;
    END
  END VDD
  OBS
      LAYER V1 ;
        RECT 0.0530 0.1010 0.0670 0.1150 ;
        RECT 0.1730 0.1010 0.1870 0.1150 ;
      LAYER V0 ;
        RECT 0.0530 0.1010 0.0670 0.1150 ;
        RECT 0.1730 0.0290 0.1870 0.0430 ;
      LAYER M0 ;
        RECT 0.0105 0.0530 0.3045 0.0670 ;
        RECT 0.0555 0.0770 0.1695 0.0910 ;
  END
END OAI21_X2

MACRO OAI21_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21_X1 0 0 ;
  SIZE 0.1800 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0430 0.0570 0.0290 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.0430 0.1575 0.0290 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0910 0.1695 0.0770 ;
    END
  END ZN
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1125 0.1010 ;
    END
  END A2
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0530 0.1245 0.0670 ;
  END
END OAI21_X1

MACRO NOR4_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4_X2 0 0 ;
  SIZE 0.4050 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0430 0.1920 0.0290 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.0430 0.3720 0.0290 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0670 0.3945 0.0530 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1470 0.1010 ;
    END
  END A1
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2580 0.1150 0.3270 0.1010 ;
    END
  END A4
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.4050 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.4050 0.1620 ;
    END
  END VDD
  OBS
      LAYER M2 ;
        RECT 0.0180 0.0290 0.3720 0.0430 ;
      LAYER V0 ;
        RECT 0.0230 0.1010 0.0370 0.1150 ;
        RECT 0.2030 0.1010 0.2170 0.1150 ;
        RECT 0.3530 0.1010 0.3670 0.1150 ;
      LAYER M1 ;
        RECT 0.0225 0.1200 0.0375 0.0240 ;
        RECT 0.2025 0.1200 0.2175 0.0240 ;
        RECT 0.3525 0.1200 0.3675 0.0240 ;
      LAYER V1 ;
        RECT 0.0230 0.0290 0.0370 0.0430 ;
        RECT 0.2030 0.0290 0.2170 0.0430 ;
        RECT 0.3530 0.0290 0.3670 0.0430 ;
      LAYER M0 ;
        RECT 0.0555 0.0770 0.1695 0.0910 ;
        RECT 0.2355 0.0770 0.3495 0.0910 ;
        RECT 0.0105 0.1010 0.0450 0.1150 ;
        RECT 0.1905 0.1010 0.2250 0.1150 ;
        RECT 0.3480 0.1010 0.3945 0.1150 ;
  END
END NOR4_X2

MACRO NOR4_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR4_X1 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0670 0.2145 0.0530 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0910 0.0570 0.0770 ;
    END
  END A1
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.0910 0.2025 0.0770 ;
    END
  END A4
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.1150 0.1020 0.1010 ;
    END
  END A2
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
END NOR4_X1

MACRO NOR3_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3_X2 0 0 ;
  SIZE 0.3150 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0180 0.0910 0.1920 0.0770 ;
      LAYER M1 ;
        RECT 0.0225 0.0960 0.0375 0.0240 ;
        RECT 0.1725 0.0960 0.1875 0.0240 ;
      LAYER M0 ;
        RECT 0.0180 0.0430 0.0570 0.0290 ;
        RECT 0.1680 0.0430 0.2025 0.0290 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.1470 0.0290 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.0670 0.2595 0.0530 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.1150 0.2820 0.1010 ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3150 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3150 0.1620 ;
    END
  END VDD
  OBS
      LAYER V1 ;
        RECT 0.0230 0.0770 0.0370 0.0910 ;
        RECT 0.1730 0.0770 0.1870 0.0910 ;
      LAYER V0 ;
        RECT 0.0230 0.0290 0.0370 0.0430 ;
        RECT 0.1730 0.0290 0.1870 0.0430 ;
      LAYER M0 ;
        RECT 0.0105 0.0770 0.3045 0.0910 ;
        RECT 0.0555 0.1010 0.1695 0.1150 ;
  END
END NOR3_X2

MACRO NOR3_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3_X1 0 0 ;
  SIZE 0.1800 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.0430 0.1020 0.0290 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0670 0.1245 0.0530 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0910 0.0570 0.0770 ;
    END
  END A1
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.1150 0.1575 0.1010 ;
    END
  END A3
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VDD
END NOR3_X1

MACRO NOR2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_X2 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0430 0.1020 0.0290 ;
    END
  END A1
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.0670 0.1695 0.0530 ;
    END
  END ZN
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.1150 0.1920 0.1010 ;
    END
  END A2
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0770 0.2145 0.0910 ;
  END
END NOR2_X2

MACRO NOR2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2_X1 0 0 ;
  SIZE 0.1350 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.1125 0.0290 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0670 0.1245 0.0530 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1150 0.0570 0.1010 ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1350 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1350 0.1620 ;
    END
  END VDD
END NOR2_X1

MACRO NAND4_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4_X2 0 0 ;
  SIZE 0.4050 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.1470 0.0290 ;
    END
  END A1
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2580 0.0430 0.3270 0.0290 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0910 0.3945 0.0770 ;
    END
  END ZN
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.1150 0.1920 0.1010 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.1150 0.3720 0.1010 ;
    END
  END A3
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.4050 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.4050 0.1620 ;
    END
  END VDD
  OBS
      LAYER M2 ;
        RECT 0.0180 0.1010 0.3720 0.1150 ;
      LAYER V0 ;
        RECT 0.0230 0.0290 0.0370 0.0430 ;
        RECT 0.2030 0.0290 0.2170 0.0430 ;
        RECT 0.3530 0.0290 0.3670 0.0430 ;
      LAYER M1 ;
        RECT 0.0225 0.1200 0.0375 0.0240 ;
        RECT 0.2025 0.1200 0.2175 0.0240 ;
        RECT 0.3525 0.1200 0.3675 0.0240 ;
      LAYER V1 ;
        RECT 0.0230 0.1010 0.0370 0.1150 ;
        RECT 0.2030 0.1010 0.2170 0.1150 ;
        RECT 0.3530 0.1010 0.3670 0.1150 ;
      LAYER M0 ;
        RECT 0.0105 0.0290 0.0450 0.0430 ;
        RECT 0.1905 0.0290 0.2250 0.0430 ;
        RECT 0.3480 0.0290 0.3945 0.0430 ;
        RECT 0.0555 0.0530 0.1695 0.0670 ;
        RECT 0.2355 0.0530 0.3495 0.0670 ;
  END
END NAND4_X2

MACRO NAND4_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND4_X1 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0670 0.0570 0.0530 ;
    END
  END A1
  PIN A4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.0670 0.2025 0.0530 ;
    END
  END A4
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0910 0.2145 0.0770 ;
    END
  END ZN
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.1150 0.1020 0.1010 ;
    END
  END A2
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
END NAND4_X1

MACRO NAND3_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3_X2 0 0 ;
  SIZE 0.3150 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0180 0.0670 0.1920 0.0530 ;
      LAYER M1 ;
        RECT 0.0225 0.1200 0.0375 0.0480 ;
        RECT 0.1725 0.1200 0.1875 0.0480 ;
      LAYER M0 ;
        RECT 0.0180 0.1150 0.0570 0.1010 ;
        RECT 0.1680 0.1150 0.2025 0.1010 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.0430 0.2820 0.0290 ;
    END
  END A1
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.0910 0.2595 0.0770 ;
    END
  END ZN
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1470 0.1010 ;
    END
  END A3
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3150 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3150 0.1620 ;
    END
  END VDD
  OBS
      LAYER V1 ;
        RECT 0.0230 0.0530 0.0370 0.0670 ;
        RECT 0.1730 0.0530 0.1870 0.0670 ;
      LAYER V0 ;
        RECT 0.0230 0.1010 0.0370 0.1150 ;
        RECT 0.1730 0.1010 0.1870 0.1150 ;
      LAYER M0 ;
        RECT 0.0555 0.0290 0.1695 0.0430 ;
        RECT 0.0105 0.0530 0.3045 0.0670 ;
  END
END NAND3_X2

MACRO NAND3_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3_X1 0 0 ;
  SIZE 0.1800 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.0430 0.1020 0.0290 ;
    END
  END A2
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0670 0.0570 0.0530 ;
    END
  END A3
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.0910 0.1695 0.0770 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.1150 0.1575 0.1010 ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VDD
END NAND3_X1

MACRO NAND2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_X2 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0430 0.1020 0.0290 ;
    END
  END A1
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.0910 0.1695 0.0770 ;
    END
  END ZN
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.1150 0.1920 0.1010 ;
    END
  END A2
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0530 0.2145 0.0670 ;
  END
END NAND2_X2

MACRO NAND2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2_X1 0 0 ;
  SIZE 0.1350 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.1125 0.0290 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0910 0.1245 0.0770 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1150 0.0570 0.1010 ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1350 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1350 0.1620 ;
    END
  END VDD
END NAND2_X1

MACRO MUX2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2_X1 0 0 ;
  SIZE 0.3150 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0430 0.1920 0.0290 ;
        RECT 0.0330 0.0910 0.1470 0.0770 ;
    END
  END S
  PIN I1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.0430 0.2475 0.0290 ;
    END
  END I1
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2700 0.0910 0.3045 0.0770 ;
    END
  END Z
  PIN I0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1125 0.1010 ;
    END
  END I0
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3150 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3150 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0530 0.1920 0.0670 ;
        RECT 0.1680 0.0770 0.2025 0.0910 ;
        RECT 0.1455 0.1010 0.2820 0.1150 ;
      LAYER V0 ;
        RECT 0.1730 0.0770 0.1870 0.0910 ;
        RECT 0.1730 0.0530 0.1870 0.0670 ;
      LAYER M1 ;
        RECT 0.1725 0.0960 0.1875 0.0240 ;
  END
END MUX2_X1

MACRO LHQ_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN LHQ_X1 0 0 ;
  SIZE 0.4500 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.3375 0.0430 0.3720 0.0290 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0670 0.0450 0.0530 ;
    END
  END Q
  PIN E
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1125 0.1010 ;
    END
  END E
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.4500 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.4500 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0330 0.0290 0.3045 0.0430 ;
        RECT 0.1005 0.0530 0.2820 0.0670 ;
        RECT 0.3030 0.0530 0.4395 0.0670 ;
        RECT 0.1005 0.0770 0.4170 0.0910 ;
        RECT 0.1455 0.1010 0.2370 0.1150 ;
        RECT 0.2580 0.1010 0.4395 0.1150 ;
  END
END LHQ_X1

MACRO INV_X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X8 0 0 ;
  SIZE 0.4050 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0430 0.3720 0.0290 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.1150 0.3495 0.1010 ;
    END
  END ZN
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.4050 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.4050 0.1620 ;
    END
  END VDD
END INV_X8

MACRO INV_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X4 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.0430 0.1695 0.0290 ;
    END
  END ZN
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.1150 0.1920 0.1010 ;
    END
  END I
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
END INV_X4

MACRO INV_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X2 0 0 ;
  SIZE 0.1350 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0430 0.1020 0.0290 ;
    END
  END I
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0450 0.1150 0.0795 0.1010 ;
    END
  END ZN
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1350 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1350 0.1620 ;
    END
  END VDD
END INV_X2

MACRO INV_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INV_X1 0 0 ;
  SIZE 0.0900 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0430 0.0795 0.0290 ;
    END
  END ZN
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1150 0.0675 0.1010 ;
    END
  END I
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.0900 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.0900 0.1620 ;
    END
  END VDD
END INV_X1

MACRO DFFRNQ_X1_SH
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFRNQ_X1_SH 0 0 ;
  SIZE 0.7650 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN RN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.3150 0.1150 0.6120 0.1010 ;
      LAYER M1 ;
        RECT 0.5925 0.1200 0.6075 0.0480 ;
        RECT 0.3225 0.1200 0.3375 0.0480 ;
      LAYER M0 ;
        RECT 0.5850 0.0670 0.6870 0.0530 ;
        RECT 0.2580 0.0670 0.3420 0.0530 ;
    END
  END RN
  PIN CK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.1150 0.0570 0.1010 ;
    END
  END CK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.7200 0.0910 0.7545 0.0770 ;
    END
  END Q
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0430 0.1125 0.0290 ;
    END
  END D
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.7650 0.1620 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.7650 0.0180 ;
    END
  END VSS
  OBS
      LAYER M2 ;
        RECT 0.1350 0.0770 0.4620 0.0910 ;
        RECT 0.1080 0.0530 0.4050 0.0670 ;
      LAYER V0 ;
        RECT 0.5930 0.0530 0.6070 0.0670 ;
        RECT 0.3230 0.0530 0.3370 0.0670 ;
        RECT 0.4430 0.0290 0.4570 0.0430 ;
        RECT 0.4430 0.1010 0.4570 0.1150 ;
        RECT 0.2030 0.0530 0.2170 0.0670 ;
        RECT 0.1430 0.1010 0.1570 0.1150 ;
        RECT 0.3830 0.0530 0.3970 0.0670 ;
        RECT 0.3830 0.1010 0.3970 0.1150 ;
        RECT 0.1130 0.0530 0.1270 0.0670 ;
        RECT 0.1130 0.0770 0.1270 0.0910 ;
      LAYER M1 ;
        RECT 0.4425 0.1200 0.4575 0.0240 ;
        RECT 0.3825 0.1200 0.3975 0.0480 ;
        RECT 0.1425 0.1200 0.1575 0.0480 ;
        RECT 0.2025 0.0960 0.2175 0.0240 ;
        RECT 0.1125 0.0960 0.1275 0.0240 ;
      LAYER V1 ;
        RECT 0.5930 0.1010 0.6070 0.1150 ;
        RECT 0.3230 0.1010 0.3370 0.1150 ;
        RECT 0.4430 0.0770 0.4570 0.0910 ;
        RECT 0.2030 0.0770 0.2170 0.0910 ;
        RECT 0.1430 0.0770 0.1570 0.0910 ;
        RECT 0.3830 0.0530 0.3970 0.0670 ;
        RECT 0.1130 0.0530 0.1270 0.0670 ;
      LAYER M0 ;
        RECT 0.6405 0.1010 0.7320 0.1150 ;
        RECT 0.4380 0.1010 0.5745 0.1150 ;
        RECT 0.3780 0.1010 0.4170 0.1150 ;
        RECT 0.1905 0.1010 0.3045 0.1150 ;
        RECT 0.1230 0.1010 0.1620 0.1150 ;
        RECT 0.4155 0.0770 0.6420 0.0910 ;
        RECT 0.2130 0.0770 0.3945 0.0910 ;
        RECT 0.1080 0.0770 0.1920 0.0910 ;
        RECT 0.3780 0.0530 0.5520 0.0670 ;
        RECT 0.1680 0.0530 0.2250 0.0670 ;
        RECT 0.0105 0.0530 0.1470 0.0670 ;
        RECT 0.4830 0.0290 0.7320 0.0430 ;
        RECT 0.3930 0.0290 0.4620 0.0430 ;
        RECT 0.1455 0.0290 0.3720 0.0430 ;
  END
END DFFRNQ_X1_SH

MACRO DFFHQN_X1_SH
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQN_X1_SH 0 0 ;
  SIZE 0.6300 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0430 0.0450 0.0290 ;
    END
  END QN
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0910 0.1125 0.0770 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.5175 0.0910 0.5520 0.0770 ;
    END
  END D
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.6300 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.6300 0.1620 ;
    END
  END VDD
  OBS
      LAYER M2 ;
        RECT 0.2880 0.0770 0.3420 0.0910 ;
      LAYER V0 ;
        RECT 0.4430 0.1010 0.4570 0.1150 ;
        RECT 0.4430 0.0530 0.4570 0.0670 ;
        RECT 0.2930 0.0770 0.3070 0.0910 ;
        RECT 0.3230 0.0290 0.3370 0.0430 ;
      LAYER M1 ;
        RECT 0.2925 0.0960 0.3075 0.0240 ;
        RECT 0.3225 0.0960 0.3375 0.0240 ;
        RECT 0.4425 0.1200 0.4575 0.0480 ;
      LAYER V1 ;
        RECT 0.2930 0.0770 0.3070 0.0910 ;
        RECT 0.3230 0.0770 0.3370 0.0910 ;
      LAYER M0 ;
        RECT 0.1005 0.0290 0.2820 0.0430 ;
        RECT 0.3030 0.0290 0.6195 0.0430 ;
        RECT 0.0330 0.0530 0.3045 0.0670 ;
        RECT 0.3255 0.0530 0.4170 0.0670 ;
        RECT 0.4380 0.0530 0.5970 0.0670 ;
        RECT 0.1455 0.0770 0.2370 0.0910 ;
        RECT 0.2580 0.0770 0.3150 0.0910 ;
        RECT 0.3480 0.0770 0.4845 0.0910 ;
        RECT 0.1005 0.1010 0.4620 0.1150 ;
        RECT 0.4830 0.1010 0.6195 0.1150 ;
  END
END DFFHQN_X1_SH

MACRO BUF_X8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X8 0 0 ;
  SIZE 0.5850 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.0430 0.1920 0.0290 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2355 0.1150 0.5295 0.1010 ;
    END
  END Z
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.5850 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.5850 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0555 0.0530 0.5520 0.0670 ;
  END
END BUF_X8

MACRO BUF_X4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X4 0 0 ;
  SIZE 0.3150 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.0430 0.2820 0.0290 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.1150 0.1695 0.1010 ;
    END
  END Z
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3150 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3150 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0330 0.0530 0.2595 0.0670 ;
  END
END BUF_X4

MACRO BUF_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X2 0 0 ;
  SIZE 0.1800 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.0430 0.1575 0.0290 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.0910 0.0900 0.0770 ;
    END
  END Z
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0330 0.1010 0.1695 0.1150 ;
  END
END BUF_X2

MACRO BUF_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUF_X1 0 0 ;
  SIZE 0.1350 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN I
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0430 0.0570 0.0290 ;
    END
  END I
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0900 0.0910 0.1245 0.0770 ;
    END
  END Z
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1350 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1350 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0105 0.1010 0.1020 0.1150 ;
  END
END BUF_X1

MACRO AOI22_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22_X2 0 0 ;
  SIZE 0.4500 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.1980 0.0670 0.2520 0.0530 ;
      LAYER M1 ;
        RECT 0.2025 0.0960 0.2175 0.0240 ;
        RECT 0.2325 0.1200 0.2475 0.0480 ;
      LAYER M0 ;
        RECT 0.1455 0.0430 0.2250 0.0290 ;
        RECT 0.2250 0.1150 0.3945 0.1010 ;
    END
  END ZN
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2580 0.0430 0.3270 0.0290 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.3480 0.0430 0.4170 0.0290 ;
    END
  END A2
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0330 0.1150 0.1020 0.1010 ;
    END
  END B2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.1150 0.1920 0.1010 ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.4500 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.4500 0.1620 ;
    END
  END VDD
  OBS
      LAYER V1 ;
        RECT 0.2030 0.0530 0.2170 0.0670 ;
        RECT 0.2330 0.0530 0.2470 0.0670 ;
      LAYER V0 ;
        RECT 0.2030 0.0290 0.2170 0.0430 ;
        RECT 0.2330 0.1010 0.2470 0.1150 ;
      LAYER M0 ;
        RECT 0.0105 0.0530 0.2145 0.0670 ;
        RECT 0.2355 0.0530 0.4395 0.0670 ;
        RECT 0.0555 0.0770 0.4395 0.0910 ;
  END
END AOI22_X2

MACRO AOI22_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22_X1 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.0525 0.1200 0.0675 0.0240 ;
      LAYER M0 ;
        RECT 0.0450 0.0430 0.1245 0.0290 ;
        RECT 0.0450 0.1150 0.0795 0.1010 ;
    END
  END ZN
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.0430 0.2025 0.0290 ;
    END
  END B2
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0670 0.0570 0.0530 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.0670 0.1125 0.0530 ;
    END
  END A1
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.1150 0.1470 0.1010 ;
    END
  END B1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  OBS
      LAYER V0 ;
        RECT 0.0530 0.1010 0.0670 0.1150 ;
        RECT 0.0530 0.0290 0.0670 0.0430 ;
      LAYER M0 ;
        RECT 0.0105 0.0770 0.2145 0.0910 ;
  END
END AOI22_X1

MACRO AOI21_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21_X2 0 0 ;
  SIZE 0.3150 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.0450 0.0670 0.1920 0.0530 ;
      LAYER M1 ;
        RECT 0.0525 0.0960 0.0675 0.0240 ;
        RECT 0.1725 0.1200 0.1875 0.0480 ;
      LAYER M0 ;
        RECT 0.0330 0.0430 0.0720 0.0290 ;
        RECT 0.1680 0.1150 0.2025 0.1010 ;
    END
  END A2
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1005 0.0430 0.2595 0.0290 ;
    END
  END ZN
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.0670 0.2820 0.0530 ;
    END
  END B
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1470 0.1010 ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.3150 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.3150 0.1620 ;
    END
  END VDD
  OBS
      LAYER V1 ;
        RECT 0.0530 0.0530 0.0670 0.0670 ;
        RECT 0.1730 0.0530 0.1870 0.0670 ;
      LAYER V0 ;
        RECT 0.0530 0.0290 0.0670 0.0430 ;
        RECT 0.1730 0.1010 0.1870 0.1150 ;
      LAYER M0 ;
        RECT 0.0555 0.0530 0.1695 0.0670 ;
        RECT 0.0105 0.0770 0.3045 0.0910 ;
  END
END AOI21_X2

MACRO AOI21_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21_X1 0 0 ;
  SIZE 0.1800 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0430 0.0570 0.0290 ;
    END
  END A1
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1230 0.0430 0.1575 0.0290 ;
    END
  END B
  PIN ZN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0105 0.0670 0.1695 0.0530 ;
    END
  END ZN
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.1150 0.1020 0.1010 ;
    END
  END A2
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0770 0.1245 0.0910 ;
  END
END AOI21_X1

MACRO AND3_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3_X2 0 0 ;
  SIZE 0.2700 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.0430 0.2025 0.0290 ;
    END
  END A3
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0555 0.0670 0.0900 0.0530 ;
    END
  END Z
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.2130 0.0670 0.2475 0.0530 ;
    END
  END A2
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.1150 0.1470 0.1010 ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2700 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2700 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0330 0.0770 0.2595 0.0910 ;
  END
END AND3_X2

MACRO AND3_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3_X1 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END A3
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0670 0.0570 0.0530 ;
    END
  END A1
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1800 0.0670 0.2145 0.0530 ;
    END
  END Z
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0780 0.1150 0.1125 0.1010 ;
    END
  END A2
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0770 0.1920 0.0910 ;
  END
END AND3_X1

MACRO AND2_X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_X2 0 0 ;
  SIZE 0.2250 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1125 0.0430 0.1470 0.0290 ;
    END
  END A2
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0450 0.1150 0.0795 0.1010 ;
    END
  END Z
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1680 0.1150 0.2025 0.1010 ;
    END
  END A1
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.2250 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.2250 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0330 0.0530 0.2145 0.0670 ;
        RECT 0.0780 0.0770 0.1695 0.0910 ;
  END
END AND2_X2

MACRO AND2_X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2_X1 0 0 ;
  SIZE 0.1800 BY 0.1440 ;
  SYMMETRY X Y ;
  SITE coresite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0225 0.0430 0.0570 0.0290 ;
    END
  END A1
  PIN Z
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.1350 0.0430 0.1695 0.0290 ;
    END
  END Z
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M0 ;
        RECT 0.0675 0.1150 0.1020 0.1010 ;
    END
  END A2
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 -0.0180 0.1800 0.0180 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M0 ;
        RECT 0.0000 0.1260 0.1800 0.1620 ;
    END
  END VDD
  OBS
      LAYER M0 ;
        RECT 0.0105 0.0530 0.1470 0.0670 ;
        RECT 0.0555 0.0770 0.1470 0.0910 ;
  END
END AND2_X1

